
module EdgeAux ( Eid, InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [11:0] Eid;
input  [11:0] WeightAddr;
input  [0:0] InEdge;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire \Weight[0] , n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, 
        n71, n72, n73, n74, n75, n76, n77;
    VMW_AND2 U15 ( .A(InEdge), .B(\Weight[0] ), .Z(OutEdge) );
    VMW_AND5 U16 ( .A(n61), .B(n62), .C(n63), .D(n64), .E(n65), .Z(n60) );
    VMW_AO22 U17 ( .A(\Weight[0] ), .B(n66), .C(WeightData), .D(n60), .Z(n77)
         );
    VMW_AND3 U18 ( .A(n68), .B(n69), .C(n70), .Z(n67) );
    VMW_AND4 U19 ( .A(n71), .B(n72), .C(n73), .D(n67), .Z(n65) );
    VMW_AND3 U20 ( .A(n74), .B(n75), .C(n76), .Z(n64) );
    VMW_XNOR2 U21 ( .A(WeightAddr[8]), .B(Eid[8]), .Z(n69) );
    VMW_XNOR2 U22 ( .A(WeightAddr[10]), .B(Eid[10]), .Z(n68) );
    VMW_XNOR2 U23 ( .A(WeightAddr[9]), .B(Eid[9]), .Z(n70) );
    VMW_XNOR2 U24 ( .A(WeightAddr[5]), .B(Eid[5]), .Z(n72) );
    VMW_XNOR2 U25 ( .A(WeightAddr[7]), .B(Eid[7]), .Z(n71) );
    VMW_XNOR2 U26 ( .A(WeightAddr[6]), .B(Eid[6]), .Z(n73) );
    VMW_XNOR2 U27 ( .A(WeightAddr[0]), .B(Eid[0]), .Z(n75) );
    VMW_XNOR2 U28 ( .A(WeightAddr[4]), .B(Eid[4]), .Z(n74) );
    VMW_XNOR2 U29 ( .A(WeightAddr[2]), .B(Eid[2]), .Z(n76) );
    VMW_XNOR2 U30 ( .A(WeightAddr[11]), .B(Eid[11]), .Z(n62) );
    VMW_XNOR2 U31 ( .A(WeightAddr[1]), .B(Eid[1]), .Z(n61) );
    VMW_XNOR2 U32 ( .A(WeightAddr[3]), .B(Eid[3]), .Z(n63) );
    VMW_INV U33 ( .A(n60), .Z(n66) );
    VMW_FD \Weight_reg[0]  ( .D(n77), .CP(Clk), .Q(\Weight[0] ) );
endmodule


module NodeAux_INDEGREE1_SOURCE1 ( Nid, InEdges, OutEdge, PathAddr, PathData, 
    Start, Clk );
input  [8:0] Nid;
input  [0:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input  Start, Clk;
    wire \path[2] , \path[0] , \OutEdge95[0] , \path[1] , n188, n189, n190, 
        n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, 
        n203, n204, n205, n206;
    tri \PathData[1] , \PathData[2] , \PathData[0] ;
    assign PathData[2] = \PathData[2] ;
    assign PathData[1] = \PathData[1] ;
    assign PathData[0] = \PathData[0] ;
    VMW_AO22 U46 ( .A(n188), .B(OutEdge), .C(n189), .D(n190), .Z(
        \OutEdge95[0] ) );
    VMW_AO21 U47 ( .A(Start), .B(\path[1] ), .C(n188), .Z(n206) );
    VMW_AO21 U48 ( .A(\path[2] ), .B(Start), .C(n188), .Z(n205) );
    VMW_AO21 U49 ( .A(Start), .B(\path[0] ), .C(n188), .Z(n204) );
    VMW_AND2 U50 ( .A(InEdges), .B(n191), .Z(n190) );
    VMW_NOR2 U51 ( .A(Start), .B(n190), .Z(n188) );
    VMW_AND3 U52 ( .A(n193), .B(n194), .C(n195), .Z(n192) );
    VMW_AND4 U53 ( .A(n197), .B(n198), .C(n199), .D(n200), .Z(n196) );
    VMW_AND4 U54 ( .A(n201), .B(n202), .C(n192), .D(n196), .Z(n203) );
    VMW_XNOR2 U55 ( .A(PathAddr[2]), .B(Nid[2]), .Z(n194) );
    VMW_XNOR2 U56 ( .A(PathAddr[0]), .B(Nid[0]), .Z(n193) );
    VMW_XNOR2 U57 ( .A(PathAddr[1]), .B(Nid[1]), .Z(n195) );
    VMW_XNOR2 U58 ( .A(PathAddr[3]), .B(Nid[3]), .Z(n202) );
    VMW_XNOR2 U59 ( .A(PathAddr[4]), .B(Nid[4]), .Z(n201) );
    VMW_XNOR2 U60 ( .A(PathAddr[5]), .B(Nid[5]), .Z(n200) );
    VMW_XNOR2 U61 ( .A(PathAddr[6]), .B(Nid[6]), .Z(n199) );
    VMW_XNOR2 U62 ( .A(PathAddr[7]), .B(Nid[7]), .Z(n198) );
    VMW_XNOR2 U63 ( .A(PathAddr[8]), .B(Nid[8]), .Z(n197) );
    VMW_INV U64 ( .A(Start), .Z(n189) );
    VMW_INV U65 ( .A(OutEdge), .Z(n191) );
    VMW_BUFIZ U66 ( .A(\path[1] ), .E(n203), .Z(\PathData[1] ) );
    VMW_BUFIZ U67 ( .A(\path[0] ), .E(n203), .Z(\PathData[0] ) );
    VMW_BUFIZ U68 ( .A(\path[2] ), .E(n203), .Z(\PathData[2] ) );
    VMW_FD \path_reg[0]  ( .D(n204), .CP(Clk), .Q(\path[0] ) );
    VMW_FD \path_reg[2]  ( .D(n205), .CP(Clk), .Q(\path[2] ) );
    VMW_FD \path_reg[1]  ( .D(n206), .CP(Clk), .Q(\path[1] ) );
    VMW_FD \OutEdge_reg[0]  ( .D(\OutEdge95[0] ), .CP(Clk), .Q(OutEdge) );
endmodule


module NodeAux_INDEGREE1_SOURCE0 ( Nid, InEdges, OutEdge, PathAddr, PathData, 
    Start, Clk );
input  [8:0] Nid;
input  [0:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input  Start, Clk;
    wire \path[2] , \path[0] , \OutEdge95[0] , \path[1] , n188, n189, n190, 
        n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, 
        n203, n204, n205, n206;
    tri \PathData[1] , \PathData[2] , \PathData[0] ;
    assign PathData[2] = \PathData[2] ;
    assign PathData[1] = \PathData[1] ;
    assign PathData[0] = \PathData[0] ;
    VMW_AO22 U46 ( .A(n188), .B(OutEdge), .C(n189), .D(n190), .Z(
        \OutEdge95[0] ) );
    VMW_AO21 U47 ( .A(Start), .B(\path[1] ), .C(n188), .Z(n206) );
    VMW_AO21 U48 ( .A(\path[2] ), .B(Start), .C(n188), .Z(n205) );
    VMW_AO21 U49 ( .A(Start), .B(\path[0] ), .C(n188), .Z(n204) );
    VMW_AND2 U50 ( .A(InEdges), .B(n191), .Z(n190) );
    VMW_NOR2 U51 ( .A(Start), .B(n190), .Z(n188) );
    VMW_AND3 U52 ( .A(n193), .B(n194), .C(n195), .Z(n192) );
    VMW_AND4 U53 ( .A(n197), .B(n198), .C(n199), .D(n200), .Z(n196) );
    VMW_AND4 U54 ( .A(n201), .B(n202), .C(n192), .D(n196), .Z(n203) );
    VMW_XNOR2 U55 ( .A(PathAddr[2]), .B(Nid[2]), .Z(n194) );
    VMW_XNOR2 U56 ( .A(PathAddr[0]), .B(Nid[0]), .Z(n193) );
    VMW_XNOR2 U57 ( .A(PathAddr[1]), .B(Nid[1]), .Z(n195) );
    VMW_XNOR2 U58 ( .A(PathAddr[3]), .B(Nid[3]), .Z(n202) );
    VMW_XNOR2 U59 ( .A(PathAddr[4]), .B(Nid[4]), .Z(n201) );
    VMW_XNOR2 U60 ( .A(PathAddr[5]), .B(Nid[5]), .Z(n200) );
    VMW_XNOR2 U61 ( .A(PathAddr[6]), .B(Nid[6]), .Z(n199) );
    VMW_XNOR2 U62 ( .A(PathAddr[7]), .B(Nid[7]), .Z(n198) );
    VMW_XNOR2 U63 ( .A(PathAddr[8]), .B(Nid[8]), .Z(n197) );
    VMW_INV U64 ( .A(Start), .Z(n189) );
    VMW_INV U65 ( .A(OutEdge), .Z(n191) );
    VMW_BUFIZ U66 ( .A(\path[1] ), .E(n203), .Z(\PathData[1] ) );
    VMW_BUFIZ U67 ( .A(\path[0] ), .E(n203), .Z(\PathData[0] ) );
    VMW_BUFIZ U68 ( .A(\path[2] ), .E(n203), .Z(\PathData[2] ) );
    VMW_FD \path_reg[0]  ( .D(n204), .CP(Clk), .Q(\path[0] ) );
    VMW_FD \path_reg[2]  ( .D(n205), .CP(Clk), .Q(\path[2] ) );
    VMW_FD \path_reg[1]  ( .D(n206), .CP(Clk), .Q(\path[1] ) );
    VMW_FD \OutEdge_reg[0]  ( .D(\OutEdge95[0] ), .CP(Clk), .Q(OutEdge) );
endmodule


module NodeAux_INDEGREE2_SOURCE0 ( Nid, InEdges, OutEdge, PathAddr, PathData, 
    Start, Clk );
input  [8:0] Nid;
input  [1:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input  Start, Clk;
    wire \path[2] , \path[0] , \OutEdge105[0] , \path[1] , n213, n214, n215, 
        n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, 
        n228, n229, n230, n231, n232, n233;
    tri \PathData[1] , \PathData[2] , \PathData[0] ;
    assign PathData[2] = \PathData[2] ;
    assign PathData[1] = \PathData[1] ;
    assign PathData[0] = \PathData[0] ;
    VMW_NOR2 U55 ( .A(Start), .B(n213), .Z(\OutEdge105[0] ) );
    VMW_AO21 U56 ( .A(Start), .B(\path[1] ), .C(n214), .Z(n233) );
    VMW_AO21 U57 ( .A(\path[2] ), .B(Start), .C(n214), .Z(n232) );
    VMW_AND3 U58 ( .A(n215), .B(n216), .C(n217), .Z(n213) );
    VMW_NAND2 U59 ( .A(InEdges[0]), .B(n215), .Z(n216) );
    VMW_AO22 U60 ( .A(n216), .B(n218), .C(\path[0] ), .D(Start), .Z(n231) );
    VMW_AND3 U61 ( .A(n220), .B(n221), .C(n222), .Z(n219) );
    VMW_AND4 U62 ( .A(n224), .B(n225), .C(n226), .D(n227), .Z(n223) );
    VMW_NAND2 U63 ( .A(InEdges[1]), .B(n215), .Z(n217) );
    VMW_AND3 U64 ( .A(n216), .B(n218), .C(n217), .Z(n214) );
    VMW_AND4 U65 ( .A(n228), .B(n229), .C(n219), .D(n223), .Z(n230) );
    VMW_XNOR2 U66 ( .A(PathAddr[2]), .B(Nid[2]), .Z(n221) );
    VMW_XNOR2 U67 ( .A(PathAddr[0]), .B(Nid[0]), .Z(n220) );
    VMW_XNOR2 U68 ( .A(PathAddr[1]), .B(Nid[1]), .Z(n222) );
    VMW_XNOR2 U69 ( .A(PathAddr[3]), .B(Nid[3]), .Z(n229) );
    VMW_XNOR2 U70 ( .A(PathAddr[4]), .B(Nid[4]), .Z(n228) );
    VMW_XNOR2 U71 ( .A(PathAddr[5]), .B(Nid[5]), .Z(n227) );
    VMW_XNOR2 U72 ( .A(PathAddr[6]), .B(Nid[6]), .Z(n226) );
    VMW_XNOR2 U73 ( .A(PathAddr[7]), .B(Nid[7]), .Z(n225) );
    VMW_XNOR2 U74 ( .A(PathAddr[8]), .B(Nid[8]), .Z(n224) );
    VMW_INV U75 ( .A(Start), .Z(n218) );
    VMW_INV U76 ( .A(OutEdge), .Z(n215) );
    VMW_BUFIZ U77 ( .A(\path[1] ), .E(n230), .Z(\PathData[1] ) );
    VMW_BUFIZ U78 ( .A(\path[0] ), .E(n230), .Z(\PathData[0] ) );
    VMW_BUFIZ U79 ( .A(\path[2] ), .E(n230), .Z(\PathData[2] ) );
    VMW_FD \path_reg[0]  ( .D(n231), .CP(Clk), .Q(\path[0] ) );
    VMW_FD \path_reg[2]  ( .D(n232), .CP(Clk), .Q(\path[2] ) );
    VMW_FD \path_reg[1]  ( .D(n233), .CP(Clk), .Q(\path[1] ) );
    VMW_FD \OutEdge_reg[0]  ( .D(\OutEdge105[0] ), .CP(Clk), .Q(OutEdge) );
endmodule


module NodeAux_INDEGREE3_SOURCE0 ( Nid, InEdges, OutEdge, PathAddr, PathData, 
    Start, Clk );
input  [8:0] Nid;
input  [2:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input  Start, Clk;
    wire \path[2] , \path[0] , \path[1] , \OutEdge115[0] , n238, n239, n240, 
        n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, 
        n253, n254, n255, n256, n257, n258, n259, n260;
    tri \PathData[1] , \PathData[2] , \PathData[0] ;
    assign PathData[2] = \PathData[2] ;
    assign PathData[1] = \PathData[1] ;
    assign PathData[0] = \PathData[0] ;
    VMW_AOI21 U64 ( .A(n238), .B(n239), .C(Start), .Z(\OutEdge115[0] ) );
    VMW_AO21 U65 ( .A(Start), .B(\path[1] ), .C(n240), .Z(n260) );
    VMW_AO22 U66 ( .A(\path[2] ), .B(Start), .C(n239), .D(n240), .Z(n259) );
    VMW_NOR3 U67 ( .A(InEdges[1]), .B(n241), .C(OutEdge), .Z(n238) );
    VMW_AOI211 U68 ( .A(n242), .B(InEdges[1]), .C(n241), .D(Start), .Z(n240)
         );
    VMW_MUX2I U69 ( .A(n243), .B(n244), .S(Start), .Z(n258) );
    VMW_AND3 U70 ( .A(n246), .B(n247), .C(n248), .Z(n245) );
    VMW_AND4 U71 ( .A(n250), .B(n251), .C(n252), .D(n253), .Z(n249) );
    VMW_NAND2 U72 ( .A(InEdges[0]), .B(n242), .Z(n254) );
    VMW_NAND2 U73 ( .A(InEdges[2]), .B(n238), .Z(n239) );
    VMW_AND4 U74 ( .A(n255), .B(n256), .C(n245), .D(n249), .Z(n257) );
    VMW_XNOR2 U75 ( .A(PathAddr[2]), .B(Nid[2]), .Z(n247) );
    VMW_XNOR2 U76 ( .A(PathAddr[0]), .B(Nid[0]), .Z(n246) );
    VMW_XNOR2 U77 ( .A(PathAddr[1]), .B(Nid[1]), .Z(n248) );
    VMW_XNOR2 U78 ( .A(PathAddr[3]), .B(Nid[3]), .Z(n256) );
    VMW_XNOR2 U79 ( .A(PathAddr[4]), .B(Nid[4]), .Z(n255) );
    VMW_XNOR2 U80 ( .A(PathAddr[5]), .B(Nid[5]), .Z(n253) );
    VMW_XNOR2 U81 ( .A(PathAddr[6]), .B(Nid[6]), .Z(n252) );
    VMW_XNOR2 U82 ( .A(PathAddr[7]), .B(Nid[7]), .Z(n251) );
    VMW_XNOR2 U83 ( .A(PathAddr[8]), .B(Nid[8]), .Z(n250) );
    VMW_NAND2 U84 ( .A(n239), .B(n254), .Z(n243) );
    VMW_INV U85 ( .A(OutEdge), .Z(n242) );
    VMW_INV U86 ( .A(\path[0] ), .Z(n244) );
    VMW_INV U87 ( .A(n254), .Z(n241) );
    VMW_BUFIZ U88 ( .A(\path[1] ), .E(n257), .Z(\PathData[1] ) );
    VMW_BUFIZ U89 ( .A(\path[0] ), .E(n257), .Z(\PathData[0] ) );
    VMW_BUFIZ U90 ( .A(\path[2] ), .E(n257), .Z(\PathData[2] ) );
    VMW_FD \path_reg[0]  ( .D(n258), .CP(Clk), .Q(\path[0] ) );
    VMW_FD \path_reg[2]  ( .D(n259), .CP(Clk), .Q(\path[2] ) );
    VMW_FD \path_reg[1]  ( .D(n260), .CP(Clk), .Q(\path[1] ) );
    VMW_FD \OutEdge_reg[0]  ( .D(\OutEdge115[0] ), .CP(Clk), .Q(OutEdge) );
endmodule


module NodeAux_INDEGREE4_SOURCE0 ( Nid, InEdges, OutEdge, PathAddr, PathData, 
    Start, Clk );
input  [8:0] Nid;
input  [3:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input  Start, Clk;
    wire \path[2] , \path[0] , \OutEdge125[0] , \path[1] , n263, n264, n265, 
        n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, 
        n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, 
        n290;
    tri \PathData[1] , \PathData[2] , \PathData[0] ;
    assign PathData[2] = \PathData[2] ;
    assign PathData[1] = \PathData[1] ;
    assign PathData[0] = \PathData[0] ;
    VMW_NOR2 U73 ( .A(Start), .B(n263), .Z(\OutEdge125[0] ) );
    VMW_AO21 U74 ( .A(n265), .B(InEdges[1]), .C(n266), .Z(n264) );
    VMW_OR3 U75 ( .A(InEdges[1]), .B(OutEdge), .C(InEdges[0]), .Z(n267) );
    VMW_NOR3 U76 ( .A(n268), .B(n269), .C(n267), .Z(n263) );
    VMW_MUX2I U77 ( .A(n270), .B(n271), .S(Start), .Z(n289) );
    VMW_MUX2I U78 ( .A(n264), .B(n272), .S(Start), .Z(n290) );
    VMW_MUX2I U79 ( .A(n273), .B(n274), .S(Start), .Z(n288) );
    VMW_AND3 U80 ( .A(n276), .B(n277), .C(n278), .Z(n275) );
    VMW_AND4 U81 ( .A(n280), .B(n281), .C(n282), .D(n283), .Z(n279) );
    VMW_AND2 U82 ( .A(n265), .B(InEdges[0]), .Z(n266) );
    VMW_AND2 U83 ( .A(InEdges[2]), .B(n284), .Z(n269) );
    VMW_AND2 U84 ( .A(InEdges[3]), .B(n284), .Z(n268) );
    VMW_AND4 U85 ( .A(n285), .B(n286), .C(n275), .D(n279), .Z(n287) );
    VMW_XNOR2 U86 ( .A(PathAddr[2]), .B(Nid[2]), .Z(n277) );
    VMW_XNOR2 U87 ( .A(PathAddr[0]), .B(Nid[0]), .Z(n276) );
    VMW_XNOR2 U88 ( .A(PathAddr[1]), .B(Nid[1]), .Z(n278) );
    VMW_XNOR2 U89 ( .A(PathAddr[3]), .B(Nid[3]), .Z(n286) );
    VMW_XNOR2 U90 ( .A(PathAddr[4]), .B(Nid[4]), .Z(n285) );
    VMW_XNOR2 U91 ( .A(PathAddr[5]), .B(Nid[5]), .Z(n283) );
    VMW_XNOR2 U92 ( .A(PathAddr[6]), .B(Nid[6]), .Z(n282) );
    VMW_XNOR2 U93 ( .A(PathAddr[7]), .B(Nid[7]), .Z(n281) );
    VMW_XNOR2 U94 ( .A(PathAddr[8]), .B(Nid[8]), .Z(n280) );
    VMW_OR3 U95 ( .A(n268), .B(n269), .C(n264), .Z(n270) );
    VMW_OR2 U96 ( .A(n266), .B(n269), .Z(n273) );
    VMW_INV U97 ( .A(OutEdge), .Z(n265) );
    VMW_INV U98 ( .A(\path[2] ), .Z(n271) );
    VMW_INV U99 ( .A(\path[0] ), .Z(n274) );
    VMW_INV U100 ( .A(\path[1] ), .Z(n272) );
    VMW_INV U101 ( .A(n267), .Z(n284) );
    VMW_BUFIZ U102 ( .A(\path[1] ), .E(n287), .Z(\PathData[1] ) );
    VMW_BUFIZ U103 ( .A(\path[0] ), .E(n287), .Z(\PathData[0] ) );
    VMW_BUFIZ U104 ( .A(\path[2] ), .E(n287), .Z(\PathData[2] ) );
    VMW_FD \path_reg[0]  ( .D(n288), .CP(Clk), .Q(\path[0] ) );
    VMW_FD \path_reg[2]  ( .D(n289), .CP(Clk), .Q(\path[2] ) );
    VMW_FD \path_reg[1]  ( .D(n290), .CP(Clk), .Q(\path[1] ) );
    VMW_FD \OutEdge_reg[0]  ( .D(\OutEdge125[0] ), .CP(Clk), .Q(OutEdge) );
endmodule


module NodeAux_INDEGREE5_SOURCE0 ( Nid, InEdges, OutEdge, PathAddr, PathData, 
    Start, Clk );
input  [8:0] Nid;
input  [4:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input  Start, Clk;
    wire \path[2] , \path[0] , \OutEdge135[0] , \path[1] , n288, n289, n290, 
        n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, 
        n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, 
        n315, n316;
    tri \PathData[1] , \PathData[2] , \PathData[0] ;
    assign PathData[2] = \PathData[2] ;
    assign PathData[1] = \PathData[1] ;
    assign PathData[0] = \PathData[0] ;
    VMW_OAI22 U82 ( .A(n288), .B(n289), .C(Start), .D(n290), .Z(
        \OutEdge135[0] ) );
    VMW_OAI22 U83 ( .A(n291), .B(n292), .C(n293), .D(n289), .Z(n316) );
    VMW_OAI22 U84 ( .A(n291), .B(n294), .C(n289), .D(n295), .Z(n314) );
    VMW_AO21 U85 ( .A(n296), .B(InEdges[1]), .C(n297), .Z(n293) );
    VMW_NOR3 U86 ( .A(InEdges[1]), .B(OutEdge), .C(InEdges[0]), .Z(n298) );
    VMW_NOR3 U87 ( .A(InEdges[2]), .B(InEdges[3]), .C(n299), .Z(n288) );
    VMW_NAND2 U88 ( .A(n291), .B(n290), .Z(n289) );
    VMW_NAND2 U89 ( .A(InEdges[4]), .B(n288), .Z(n290) );
    VMW_AO22 U90 ( .A(n300), .B(n291), .C(\path[2] ), .D(Start), .Z(n315) );
    VMW_OR2 U91 ( .A(n297), .B(n301), .Z(n295) );
    VMW_AND3 U92 ( .A(n303), .B(n304), .C(n305), .Z(n302) );
    VMW_AND4 U93 ( .A(n307), .B(n308), .C(n309), .D(n310), .Z(n306) );
    VMW_AND2 U94 ( .A(n296), .B(InEdges[0]), .Z(n297) );
    VMW_AND2 U95 ( .A(n298), .B(InEdges[2]), .Z(n301) );
    VMW_AND4 U96 ( .A(n311), .B(n312), .C(n302), .D(n306), .Z(n313) );
    VMW_XNOR2 U97 ( .A(PathAddr[2]), .B(Nid[2]), .Z(n304) );
    VMW_XNOR2 U98 ( .A(PathAddr[0]), .B(Nid[0]), .Z(n303) );
    VMW_XNOR2 U99 ( .A(PathAddr[1]), .B(Nid[1]), .Z(n305) );
    VMW_XNOR2 U100 ( .A(PathAddr[3]), .B(Nid[3]), .Z(n312) );
    VMW_XNOR2 U101 ( .A(PathAddr[4]), .B(Nid[4]), .Z(n311) );
    VMW_XNOR2 U102 ( .A(PathAddr[5]), .B(Nid[5]), .Z(n310) );
    VMW_XNOR2 U103 ( .A(PathAddr[6]), .B(Nid[6]), .Z(n309) );
    VMW_XNOR2 U104 ( .A(PathAddr[7]), .B(Nid[7]), .Z(n308) );
    VMW_XNOR2 U105 ( .A(PathAddr[8]), .B(Nid[8]), .Z(n307) );
    VMW_AOI211 U106 ( .A(n298), .B(InEdges[3]), .C(n301), .D(n293), .Z(n300)
         );
    VMW_INV U107 ( .A(Start), .Z(n291) );
    VMW_INV U108 ( .A(OutEdge), .Z(n296) );
    VMW_INV U109 ( .A(\path[0] ), .Z(n294) );
    VMW_INV U110 ( .A(\path[1] ), .Z(n292) );
    VMW_INV U111 ( .A(n298), .Z(n299) );
    VMW_BUFIZ U112 ( .A(\path[1] ), .E(n313), .Z(\PathData[1] ) );
    VMW_BUFIZ U113 ( .A(\path[0] ), .E(n313), .Z(\PathData[0] ) );
    VMW_BUFIZ U114 ( .A(\path[2] ), .E(n313), .Z(\PathData[2] ) );
    VMW_FD \path_reg[0]  ( .D(n314), .CP(Clk), .Q(\path[0] ) );
    VMW_FD \path_reg[2]  ( .D(n315), .CP(Clk), .Q(\path[2] ) );
    VMW_FD \path_reg[1]  ( .D(n316), .CP(Clk), .Q(\path[1] ) );
    VMW_FD \OutEdge_reg[0]  ( .D(\OutEdge135[0] ), .CP(Clk), .Q(OutEdge) );
endmodule


module NodeAux_INDEGREE6_SOURCE0 ( Nid, InEdges, OutEdge, PathAddr, PathData, 
    Start, Clk );
input  [8:0] Nid;
input  [5:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input  Start, Clk;
    wire \OutEdge145[0] , \path[2] , \path[0] , \path[1] , n313, n314, n315, 
        n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, 
        n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, 
        n340, n341, n342, n343, n344;
    tri \PathData[1] , \PathData[2] , \PathData[0] ;
    assign PathData[2] = \PathData[2] ;
    assign PathData[1] = \PathData[1] ;
    assign PathData[0] = \PathData[0] ;
    VMW_NOR2 U91 ( .A(Start), .B(n313), .Z(\OutEdge145[0] ) );
    VMW_AO21 U92 ( .A(n315), .B(InEdges[1]), .C(n316), .Z(n314) );
    VMW_NOR3 U93 ( .A(InEdges[1]), .B(OutEdge), .C(InEdges[0]), .Z(n317) );
    VMW_NOR3 U94 ( .A(InEdges[2]), .B(InEdges[3]), .C(n319), .Z(n318) );
    VMW_NOR3 U95 ( .A(n320), .B(n321), .C(n322), .Z(n313) );
    VMW_AO22 U96 ( .A(n323), .B(n324), .C(\path[2] ), .D(Start), .Z(n343) );
    VMW_OAI22 U97 ( .A(n326), .B(Start), .C(\path[1] ), .D(n324), .Z(n325) );
    VMW_OAI22 U98 ( .A(n328), .B(Start), .C(\path[0] ), .D(n324), .Z(n327) );
    VMW_AND3 U99 ( .A(n330), .B(n331), .C(n332), .Z(n329) );
    VMW_AND4 U100 ( .A(n334), .B(n335), .C(n336), .D(n337), .Z(n333) );
    VMW_AND2 U101 ( .A(n315), .B(InEdges[0]), .Z(n316) );
    VMW_AND2 U102 ( .A(n317), .B(InEdges[2]), .Z(n338) );
    VMW_AND2 U103 ( .A(InEdges[4]), .B(n318), .Z(n321) );
    VMW_AND2 U104 ( .A(InEdges[5]), .B(n318), .Z(n322) );
    VMW_AND4 U105 ( .A(n339), .B(n340), .C(n329), .D(n333), .Z(n341) );
    VMW_XNOR2 U106 ( .A(PathAddr[2]), .B(Nid[2]), .Z(n331) );
    VMW_XNOR2 U107 ( .A(PathAddr[0]), .B(Nid[0]), .Z(n330) );
    VMW_XNOR2 U108 ( .A(PathAddr[1]), .B(Nid[1]), .Z(n332) );
    VMW_XNOR2 U109 ( .A(PathAddr[3]), .B(Nid[3]), .Z(n340) );
    VMW_XNOR2 U110 ( .A(PathAddr[4]), .B(Nid[4]), .Z(n339) );
    VMW_XNOR2 U111 ( .A(PathAddr[5]), .B(Nid[5]), .Z(n337) );
    VMW_XNOR2 U112 ( .A(PathAddr[6]), .B(Nid[6]), .Z(n336) );
    VMW_XNOR2 U113 ( .A(PathAddr[7]), .B(Nid[7]), .Z(n335) );
    VMW_XNOR2 U114 ( .A(PathAddr[8]), .B(Nid[8]), .Z(n334) );
    VMW_AOI211 U115 ( .A(n317), .B(InEdges[3]), .C(n338), .D(n314), .Z(n323)
         );
    VMW_NOR3 U116 ( .A(n322), .B(n321), .C(n314), .Z(n326) );
    VMW_NOR3 U117 ( .A(n338), .B(n316), .C(n321), .Z(n328) );
    VMW_INV U118 ( .A(Start), .Z(n324) );
    VMW_INV U119 ( .A(OutEdge), .Z(n315) );
    VMW_INV U120 ( .A(n317), .Z(n319) );
    VMW_INV U121 ( .A(n318), .Z(n320) );
    VMW_INV U122 ( .A(n325), .Z(n344) );
    VMW_INV U123 ( .A(n327), .Z(n342) );
    VMW_BUFIZ U124 ( .A(\path[1] ), .E(n341), .Z(\PathData[1] ) );
    VMW_BUFIZ U125 ( .A(\path[0] ), .E(n341), .Z(\PathData[0] ) );
    VMW_BUFIZ U126 ( .A(\path[2] ), .E(n341), .Z(\PathData[2] ) );
    VMW_FD \path_reg[0]  ( .D(n342), .CP(Clk), .Q(\path[0] ) );
    VMW_FD \path_reg[2]  ( .D(n343), .CP(Clk), .Q(\path[2] ) );
    VMW_FD \path_reg[1]  ( .D(n344), .CP(Clk), .Q(\path[1] ) );
    VMW_FD \OutEdge_reg[0]  ( .D(\OutEdge145[0] ), .CP(Clk), .Q(OutEdge) );
endmodule


module NodeAux_INDEGREE7_SOURCE0 ( Nid, InEdges, OutEdge, PathAddr, PathData, 
    Start, Clk );
input  [8:0] Nid;
input  [6:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input  Start, Clk;
    wire \path[2] , \path[0] , \path[1] , \OutEdge155[0] , n338, n339, n340, 
        n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, 
        n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, 
        n365, n366, n367, n368, n369, n370, n371, n372;
    tri \PathData[1] , \PathData[2] , \PathData[0] ;
    assign PathData[2] = \PathData[2] ;
    assign PathData[1] = \PathData[1] ;
    assign PathData[0] = \PathData[0] ;
    VMW_AOI21 U100 ( .A(n338), .B(n339), .C(Start), .Z(\OutEdge155[0] ) );
    VMW_AOI21 U101 ( .A(n341), .B(InEdges[1]), .C(n342), .Z(n340) );
    VMW_OR3 U102 ( .A(OutEdge), .B(n342), .C(InEdges[1]), .Z(n343) );
    VMW_NOR3 U103 ( .A(InEdges[2]), .B(InEdges[3]), .C(n343), .Z(n344) );
    VMW_NOR3 U104 ( .A(InEdges[5]), .B(InEdges[4]), .C(n345), .Z(n338) );
    VMW_MUX2I U105 ( .A(n346), .B(n347), .S(Start), .Z(n371) );
    VMW_MUX2I U106 ( .A(n348), .B(n349), .S(Start), .Z(n372) );
    VMW_MUX2I U107 ( .A(n350), .B(n351), .S(Start), .Z(n370) );
    VMW_AND3 U108 ( .A(n353), .B(n354), .C(n355), .Z(n352) );
    VMW_AND4 U109 ( .A(n357), .B(n358), .C(n359), .D(n360), .Z(n356) );
    VMW_NAND2 U110 ( .A(InEdges[0]), .B(n341), .Z(n361) );
    VMW_OR2 U111 ( .A(n363), .B(n343), .Z(n362) );
    VMW_NAND2 U112 ( .A(InEdges[4]), .B(n344), .Z(n364) );
    VMW_NAND2 U113 ( .A(InEdges[6]), .B(n338), .Z(n339) );
    VMW_AND4 U114 ( .A(n365), .B(n366), .C(n352), .D(n356), .Z(n369) );
    VMW_XNOR2 U115 ( .A(PathAddr[2]), .B(Nid[2]), .Z(n354) );
    VMW_XNOR2 U116 ( .A(PathAddr[0]), .B(Nid[0]), .Z(n353) );
    VMW_XNOR2 U117 ( .A(PathAddr[1]), .B(Nid[1]), .Z(n355) );
    VMW_XNOR2 U118 ( .A(PathAddr[3]), .B(Nid[3]), .Z(n366) );
    VMW_XNOR2 U119 ( .A(PathAddr[4]), .B(Nid[4]), .Z(n365) );
    VMW_XNOR2 U120 ( .A(PathAddr[5]), .B(Nid[5]), .Z(n360) );
    VMW_XNOR2 U121 ( .A(PathAddr[6]), .B(Nid[6]), .Z(n359) );
    VMW_XNOR2 U122 ( .A(PathAddr[7]), .B(Nid[7]), .Z(n358) );
    VMW_XNOR2 U123 ( .A(PathAddr[8]), .B(Nid[8]), .Z(n357) );
    VMW_OAI211 U124 ( .A(n343), .B(n367), .C(n362), .D(n340), .Z(n346) );
    VMW_OAI211 U125 ( .A(n345), .B(n368), .C(n364), .D(n340), .Z(n348) );
    VMW_NAND4 U126 ( .A(n339), .B(n364), .C(n362), .D(n361), .Z(n350) );
    VMW_INV U127 ( .A(OutEdge), .Z(n341) );
    VMW_INV U128 ( .A(InEdges[3]), .Z(n367) );
    VMW_INV U129 ( .A(n361), .Z(n342) );
    VMW_INV U130 ( .A(InEdges[5]), .Z(n368) );
    VMW_INV U131 ( .A(\path[2] ), .Z(n347) );
    VMW_INV U132 ( .A(\path[0] ), .Z(n351) );
    VMW_INV U133 ( .A(\path[1] ), .Z(n349) );
    VMW_INV U134 ( .A(InEdges[2]), .Z(n363) );
    VMW_INV U135 ( .A(n344), .Z(n345) );
    VMW_BUFIZ U136 ( .A(\path[1] ), .E(n369), .Z(\PathData[1] ) );
    VMW_BUFIZ U137 ( .A(\path[0] ), .E(n369), .Z(\PathData[0] ) );
    VMW_BUFIZ U138 ( .A(\path[2] ), .E(n369), .Z(\PathData[2] ) );
    VMW_FD \path_reg[0]  ( .D(n370), .CP(Clk), .Q(\path[0] ) );
    VMW_FD \path_reg[2]  ( .D(n371), .CP(Clk), .Q(\path[2] ) );
    VMW_FD \path_reg[1]  ( .D(n372), .CP(Clk), .Q(\path[1] ) );
    VMW_FD \OutEdge_reg[0]  ( .D(\OutEdge155[0] ), .CP(Clk), .Q(OutEdge) );
endmodule


module library ( InEdges, OutEdge, PathAddr, PathData, WeightAddr, WeightData, 
    Nid, Eid, Start, Clk );
input  [6:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
input  [11:0] WeightAddr;
input  [11:0] Eid;
output [2:0] PathData;
input  [0:0] WeightData;
input  [8:0] Nid;
input  Start, Clk;
    EdgeAux edgeAux ( .Eid(Eid), .InEdge(InEdges[0]), .OutEdge(OutEdge), 
        .WeightAddr(WeightAddr), .WeightData(WeightData), .Clk(Clk) );
    NodeAux_INDEGREE1_SOURCE1 n_1_1 ( .Nid(Nid), .InEdges(InEdges[0]), 
        .OutEdge(OutEdge), .PathAddr(PathAddr), .PathData(PathData), .Start(
        Start), .Clk(Clk) );
    NodeAux_INDEGREE1_SOURCE0 n_1_0 ( .Nid(Nid), .InEdges(InEdges[0]), 
        .OutEdge(OutEdge), .PathAddr(PathAddr), .PathData(PathData), .Start(
        Start), .Clk(Clk) );
    NodeAux_INDEGREE4_SOURCE0 n_4_0 ( .Nid(Nid), .InEdges(InEdges[3:0]), 
        .OutEdge(OutEdge), .PathAddr(PathAddr), .PathData(PathData), .Start(
        Start), .Clk(Clk) );
    NodeAux_INDEGREE5_SOURCE0 n_5_0 ( .Nid(Nid), .InEdges(InEdges[4:0]), 
        .OutEdge(OutEdge), .PathAddr(PathAddr), .PathData(PathData), .Start(
        Start), .Clk(Clk) );
    NodeAux_INDEGREE2_SOURCE0 n_2_0 ( .Nid(Nid), .InEdges(InEdges[1:0]), 
        .OutEdge(OutEdge), .PathAddr(PathAddr), .PathData(PathData), .Start(
        Start), .Clk(Clk) );
    NodeAux_INDEGREE6_SOURCE0 n_6_0 ( .Nid(Nid), .InEdges(InEdges[5:0]), 
        .OutEdge(OutEdge), .PathAddr(PathAddr), .PathData(PathData), .Start(
        Start), .Clk(Clk) );
    NodeAux_INDEGREE7_SOURCE0 n_7_0 ( .Nid(Nid), .InEdges(InEdges), .OutEdge(
        OutEdge), .PathAddr(PathAddr), .PathData(PathData), .Start(Start), 
        .Clk(Clk) );
    NodeAux_INDEGREE3_SOURCE0 n_3_0 ( .Nid(Nid), .InEdges(InEdges[2:0]), 
        .OutEdge(OutEdge), .PathAddr(PathAddr), .PathData(PathData), .Start(
        Start), .Clk(Clk) );
endmodule



module Node_NID0_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [0:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE1 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid0 , nid0 , nid0 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID0 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID1_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [5:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid0 , nid0 , nid0 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID2 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID3 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID4 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID5 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID6 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID2_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [3:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid0 , nid0 , nid0 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID7 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID8 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID9 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID10 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID3_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [5:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid0 , nid0 , nid0 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID11 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID12 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID13 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID14 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID15 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID16 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID4_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [6:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid0 , nid0 , nid0 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID17 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID18 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID19 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID20 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID21 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID22 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID23 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID5_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [0:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid0 , nid0 , nid0 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID24 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID6_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [6:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid0 , nid0 , nid0 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID25 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID26 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID27 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID28 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID29 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID30 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID31 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID7_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [3:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid0 , nid0 , nid0 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID32 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID33 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID34 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID35 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID8_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [6:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid0 , nid0 , nid1 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID36 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID37 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID38 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID39 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID40 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID41 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID42 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID9_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [5:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid0 , nid0 , nid1 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID43 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID44 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID45 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID46 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID47 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID48 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID10_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [5:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid0 , nid0 , nid1 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID49 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID50 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID51 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID52 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID53 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID54 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID11_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [3:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid0 , nid0 , nid1 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID55 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID56 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID57 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID58 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID12_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [5:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid0 , nid0 , nid1 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID59 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID60 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID61 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID62 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID63 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID64 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID13_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [5:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid0 , nid0 , nid1 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID65 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID66 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID67 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID68 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID69 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID70 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID14_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [4:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid0 , nid0 , nid1 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID71 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID72 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID73 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID74 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID75 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID15_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [1:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid0 , nid0 , nid1 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID76 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID77 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID16_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [3:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid0 , nid1 , nid0 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID78 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID79 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID80 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID81 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID17_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [1:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid0 , nid1 , nid0 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID82 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID83 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID18_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [5:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid0 , nid1 , nid0 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID84 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID85 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID86 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID87 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID88 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID89 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID19_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [6:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid0 , nid1 , nid0 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID90 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID91 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID92 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID93 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID94 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID95 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID96 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID20_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [6:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid0 , nid1 , nid0 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID97 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID98 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID99 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID100 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID101 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID102 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID103 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID21_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [3:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid0 , nid1 , nid0 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID104 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID105 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID106 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID107 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID22_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [6:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid0 , nid1 , nid0 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID108 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID109 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID110 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID111 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID112 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID113 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID114 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID23_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [3:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid0 , nid1 , nid0 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID115 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID116 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID117 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID118 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID24_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [0:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid0 , nid1 , nid1 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID119 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID25_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [6:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid0 , nid1 , nid1 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID120 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID121 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID122 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID123 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID124 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID125 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID126 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID26_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [4:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid0 , nid1 , nid1 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID127 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID128 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID129 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID130 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID131 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID27_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [5:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid0 , nid1 , nid1 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID132 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID133 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID134 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID135 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID136 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID137 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID28_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [0:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid0 , nid1 , nid1 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID138 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID29_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [2:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid0 , nid1 , nid1 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID139 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID140 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID141 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID30_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [0:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid0 , nid1 , nid1 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID142 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID31_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [5:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid0 , nid1 , nid1 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID143 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID144 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID145 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID146 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID147 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID148 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID32_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [1:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid1 , nid0 , nid0 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID149 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID150 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID33_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [6:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid1 , nid0 , nid0 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID151 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID152 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID153 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID154 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID155 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID156 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID157 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID34_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [2:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid1 , nid0 , nid0 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID158 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID159 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID160 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID35_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [5:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid1 , nid0 , nid0 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID161 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID162 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID163 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID164 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID165 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID166 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID36_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [4:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid1 , nid0 , nid0 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID167 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID168 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID169 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID170 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID171 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID37_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [6:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid1 , nid0 , nid0 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID172 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID173 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID174 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID175 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID176 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID177 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID178 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID38_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [5:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid1 , nid0 , nid0 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID179 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID180 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID181 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID182 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID183 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID184 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID39_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [1:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid1 , nid0 , nid0 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID185 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID186 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID40_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [4:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid1 , nid0 , nid1 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID187 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID188 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID189 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID190 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID191 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID41_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [0:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid1 , nid0 , nid1 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID192 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID42_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [4:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid1 , nid0 , nid1 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID193 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID194 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID195 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID196 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID197 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID43_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [2:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid1 , nid0 , nid1 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID198 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID199 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID200 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID44_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [0:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid1 , nid0 , nid1 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID201 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID45_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [2:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid1 , nid0 , nid1 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID202 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID203 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID204 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID46_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [2:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid1 , nid0 , nid1 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID205 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID206 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID207 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID47_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [3:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid1 , nid0 , nid1 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID208 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID209 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID210 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID211 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID48_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [0:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid1 , nid1 , nid0 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID212 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID49_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [6:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid1 , nid1 , nid0 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID213 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID214 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID215 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID216 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID217 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID218 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID219 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID50_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [4:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid1 , nid1 , nid0 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID220 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID221 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID222 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID223 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID224 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID51_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [6:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid1 , nid1 , nid0 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID225 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID226 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID227 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID228 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID229 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID230 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID231 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID52_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [3:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid1 , nid1 , nid0 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID232 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID233 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID234 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID235 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID53_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [0:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid1 , nid1 , nid0 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID236 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID54_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [0:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid1 , nid1 , nid0 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID237 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID55_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [4:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid1 , nid1 , nid0 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID238 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID239 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID240 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID241 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID242 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID56_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [4:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid1 , nid1 , nid1 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID243 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID244 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID245 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID246 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID247 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID57_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [2:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid1 , nid1 , nid1 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID248 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID249 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID250 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID58_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [5:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid1 , nid1 , nid1 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID251 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID252 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID253 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID254 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID255 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID256 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID59_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [2:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid1 , nid1 , nid1 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID257 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID258 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID259 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID60_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [2:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid1 , nid1 , nid1 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID260 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID261 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID262 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID61_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [0:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid1 , nid1 , nid1 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID263 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID62_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [4:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid1 , nid1 , nid1 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID264 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID265 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID266 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID267 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID268 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID63_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [4:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid0 , nid1 , nid1 , nid1 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID269 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID270 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID271 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID272 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID273 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID64_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [1:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid0 , nid0 , nid0 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID274 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID275 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID65_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [4:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid0 , nid0 , nid0 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID276 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID277 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID278 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID279 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID280 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID66_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [4:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid0 , nid0 , nid0 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID281 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID282 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID283 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID284 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID285 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID67_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [1:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid0 , nid0 , nid0 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID286 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID287 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID68_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [4:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid0 , nid0 , nid0 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID288 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID289 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID290 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID291 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID292 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID69_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [3:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid0 , nid0 , nid0 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID293 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID294 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID295 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID296 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID70_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [0:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid0 , nid0 , nid0 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID297 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID71_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [3:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid0 , nid0 , nid0 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID298 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID299 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID300 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID301 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID72_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [6:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid0 , nid0 , nid1 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID302 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID303 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID304 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID305 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID306 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID307 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID308 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID73_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [0:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid0 , nid0 , nid1 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID309 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID74_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [4:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid0 , nid0 , nid1 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID310 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID311 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID312 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID313 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID314 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID75_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [1:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid0 , nid0 , nid1 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID315 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID316 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID76_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [2:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid0 , nid0 , nid1 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID317 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID318 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID319 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID77_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [4:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid0 , nid0 , nid1 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID320 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID321 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID322 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID323 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID324 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID78_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [6:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid0 , nid0 , nid1 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID325 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID326 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID327 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID328 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID329 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID330 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID331 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID79_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [2:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid0 , nid0 , nid1 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID332 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID333 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID334 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID80_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [6:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid0 , nid1 , nid0 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID335 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID336 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID337 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID338 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID339 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID340 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID341 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID81_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [0:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid0 , nid1 , nid0 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID342 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID82_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [0:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid0 , nid1 , nid0 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID343 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID83_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [5:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid0 , nid1 , nid0 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID344 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID345 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID346 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID347 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID348 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID349 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID84_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [4:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid0 , nid1 , nid0 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID350 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID351 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID352 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID353 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID354 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID85_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [1:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid0 , nid1 , nid0 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID355 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID356 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID86_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [0:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid0 , nid1 , nid0 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID357 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID87_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [2:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid0 , nid1 , nid0 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID358 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID359 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID360 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID88_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [4:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid0 , nid1 , nid1 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID361 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID362 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID363 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID364 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID365 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID89_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [6:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid0 , nid1 , nid1 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID366 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID367 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID368 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID369 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID370 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID371 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID372 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID90_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [2:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid0 , nid1 , nid1 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID373 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID374 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID375 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID91_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [5:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid0 , nid1 , nid1 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID376 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID377 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID378 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID379 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID380 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID381 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID92_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [5:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid0 , nid1 , nid1 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID382 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID383 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID384 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID385 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID386 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID387 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID93_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [2:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid0 , nid1 , nid1 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID388 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID389 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID390 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID94_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [0:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid0 , nid1 , nid1 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID391 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID95_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [5:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid0 , nid1 , nid1 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID392 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID393 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID394 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID395 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID396 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID397 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID96_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [4:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid1 , nid0 , nid0 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID398 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID399 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID400 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID401 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID402 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID97_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [3:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid1 , nid0 , nid0 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID403 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID404 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID405 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID406 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID98_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [5:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid1 , nid0 , nid0 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID407 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID408 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID409 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID410 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID411 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID412 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID99_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [4:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid1 , nid0 , nid0 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID413 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID414 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID415 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID416 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID417 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID100_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [3:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid1 , nid0 , nid0 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID418 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID419 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID420 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID421 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID101_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [3:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid1 , nid0 , nid0 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID422 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID423 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID424 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID425 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID102_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [3:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid1 , nid0 , nid0 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID426 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID427 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID428 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID429 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID103_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [2:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid1 , nid0 , nid0 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID430 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID431 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID432 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID104_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [4:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid1 , nid0 , nid1 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID433 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID434 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID435 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID436 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID437 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID105_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [2:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid1 , nid0 , nid1 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID438 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID439 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID440 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID106_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [6:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid1 , nid0 , nid1 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID441 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID442 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID443 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID444 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID445 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID446 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID447 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID107_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [4:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid1 , nid0 , nid1 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID448 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID449 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID450 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID451 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID452 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID108_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [4:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid1 , nid0 , nid1 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID453 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID454 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID455 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID456 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID457 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID109_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [1:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid1 , nid0 , nid1 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID458 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID459 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID110_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [4:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid1 , nid0 , nid1 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID460 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID461 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID462 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID463 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID464 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID111_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [6:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid1 , nid0 , nid1 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID465 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID466 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID467 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID468 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID469 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID470 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID471 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID112_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [4:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid1 , nid1 , nid0 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID472 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID473 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID474 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID475 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID476 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID113_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [1:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid1 , nid1 , nid0 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID477 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID478 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID114_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [2:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid1 , nid1 , nid0 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID479 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID480 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID481 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID115_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [3:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid1 , nid1 , nid0 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID482 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID483 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID484 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID485 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID116_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [6:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid1 , nid1 , nid0 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID486 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID487 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID488 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID489 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID490 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID491 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID492 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID117_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [1:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid1 , nid1 , nid0 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID493 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID494 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID118_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [1:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid1 , nid1 , nid0 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID495 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID496 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID119_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [6:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid1 , nid1 , nid0 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID497 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID498 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID499 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID500 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID501 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID502 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID503 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID120_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [5:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid1 , nid1 , nid1 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID504 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID505 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID506 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID507 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID508 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID509 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID121_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [5:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid1 , nid1 , nid1 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID510 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID511 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID512 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID513 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID514 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID515 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID122_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [6:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid1 , nid1 , nid1 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID516 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID517 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID518 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID519 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID520 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID521 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID522 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID123_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [0:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid1 , nid1 , nid1 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID523 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID124_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [2:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid1 , nid1 , nid1 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID524 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID525 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID526 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID125_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [0:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid1 , nid1 , nid1 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID527 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID126_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [4:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid1 , nid1 , nid1 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID528 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID529 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID530 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID531 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID532 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID127_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [5:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid0 , nid0 , nid1 , nid1 , nid1 , nid1 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID533 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID534 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID535 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID536 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID537 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID538 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID128_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [2:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid0 , nid0 , nid0 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID539 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID540 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID541 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID129_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [2:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid0 , nid0 , nid0 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID542 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID543 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID544 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID130_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [1:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid0 , nid0 , nid0 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID545 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID546 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID131_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [3:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid0 , nid0 , nid0 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID547 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID548 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID549 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID550 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID132_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [4:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid0 , nid0 , nid0 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID551 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID552 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID553 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID554 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID555 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID133_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [6:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid0 , nid0 , nid0 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID556 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID557 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID558 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID559 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID560 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID561 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID562 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID134_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [2:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid0 , nid0 , nid0 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID563 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID564 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID565 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID135_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [6:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid0 , nid0 , nid0 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID566 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID567 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID568 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID569 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID570 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID571 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID572 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID136_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [4:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid0 , nid0 , nid1 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID573 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID574 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID575 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID576 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID577 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID137_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [2:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid0 , nid0 , nid1 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID578 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID579 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID580 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID138_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [0:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid0 , nid0 , nid1 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID581 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID139_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [1:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid0 , nid0 , nid1 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID582 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID583 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID140_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [3:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid0 , nid0 , nid1 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID584 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID585 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID586 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID587 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID141_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [6:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid0 , nid0 , nid1 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID588 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID589 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID590 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID591 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID592 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID593 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID594 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID142_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [0:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid0 , nid0 , nid1 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID595 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID143_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [5:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid0 , nid0 , nid1 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID596 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID597 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID598 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID599 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID600 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID601 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID144_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [5:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid0 , nid1 , nid0 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID602 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID603 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID604 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID605 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID606 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID607 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID145_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [2:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid0 , nid1 , nid0 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID608 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID609 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID610 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID146_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [2:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid0 , nid1 , nid0 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID611 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID612 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID613 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID147_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [4:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid0 , nid1 , nid0 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID614 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID615 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID616 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID617 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID618 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID148_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [6:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid0 , nid1 , nid0 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID619 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID620 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID621 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID622 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID623 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID624 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID625 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID149_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [3:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid0 , nid1 , nid0 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID626 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID627 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID628 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID629 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID150_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [5:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid0 , nid1 , nid0 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID630 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID631 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID632 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID633 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID634 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID635 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID151_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [2:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid0 , nid1 , nid0 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID636 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID637 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID638 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID152_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [6:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid0 , nid1 , nid1 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID639 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID640 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID641 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID642 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID643 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID644 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID645 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID153_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [3:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid0 , nid1 , nid1 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID646 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID647 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID648 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID649 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID154_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [6:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid0 , nid1 , nid1 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID650 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID651 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID652 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID653 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID654 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID655 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID656 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID155_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [0:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid0 , nid1 , nid1 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID657 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID156_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [4:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid0 , nid1 , nid1 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID658 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID659 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID660 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID661 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID662 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID157_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [6:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid0 , nid1 , nid1 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID663 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID664 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID665 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID666 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID667 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID668 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID669 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID158_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [1:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid0 , nid1 , nid1 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID670 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID671 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID159_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [6:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid0 , nid1 , nid1 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID672 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID673 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID674 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID675 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID676 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID677 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID678 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID160_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [6:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid1 , nid0 , nid0 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID679 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID680 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID681 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID682 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID683 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID684 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID685 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID161_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [3:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid1 , nid0 , nid0 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID686 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID687 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID688 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID689 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID162_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [1:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid1 , nid0 , nid0 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID690 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID691 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID163_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [6:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid1 , nid0 , nid0 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID692 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID693 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID694 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID695 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID696 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID697 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID698 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID164_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [4:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid1 , nid0 , nid0 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID699 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID700 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID701 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID702 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID703 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID165_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [0:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid1 , nid0 , nid0 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID704 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID166_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [0:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid1 , nid0 , nid0 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID705 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID167_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [5:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid1 , nid0 , nid0 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID706 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID707 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID708 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID709 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID710 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID711 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID168_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [0:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid1 , nid0 , nid1 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID712 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID169_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [3:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid1 , nid0 , nid1 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID713 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID714 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID715 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID716 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID170_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [4:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid1 , nid0 , nid1 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID717 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID718 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID719 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID720 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID721 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID171_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [4:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid1 , nid0 , nid1 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID722 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID723 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID724 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID725 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID726 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID172_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [6:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid1 , nid0 , nid1 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID727 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID728 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID729 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID730 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID731 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID732 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID733 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID173_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [1:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid1 , nid0 , nid1 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID734 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID735 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID174_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [1:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid1 , nid0 , nid1 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID736 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID737 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID175_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [0:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid1 , nid0 , nid1 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID738 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID176_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [4:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid1 , nid1 , nid0 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID739 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID740 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID741 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID742 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID743 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID177_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [0:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid1 , nid1 , nid0 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID744 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID178_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [4:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid1 , nid1 , nid0 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID745 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID746 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID747 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID748 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID749 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID179_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [6:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid1 , nid1 , nid0 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID750 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID751 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID752 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID753 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID754 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID755 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID756 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID180_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [5:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid1 , nid1 , nid0 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID757 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID758 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID759 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID760 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID761 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID762 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID181_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [6:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid1 , nid1 , nid0 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID763 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID764 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID765 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID766 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID767 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID768 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID769 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID182_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [6:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid1 , nid1 , nid0 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID770 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID771 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID772 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID773 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID774 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID775 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID776 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID183_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [3:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid1 , nid1 , nid0 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID777 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID778 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID779 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID780 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID184_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [6:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid1 , nid1 , nid1 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID781 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID782 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID783 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID784 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID785 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID786 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID787 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID185_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [0:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid1 , nid1 , nid1 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID788 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID186_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [0:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid1 , nid1 , nid1 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID789 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID187_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [2:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid1 , nid1 , nid1 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID790 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID791 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID792 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID188_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [4:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid1 , nid1 , nid1 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID793 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID794 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID795 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID796 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID797 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID189_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [6:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid1 , nid1 , nid1 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID798 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID799 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID800 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID801 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID802 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID803 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID804 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID190_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [6:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid1 , nid1 , nid1 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID805 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID806 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID807 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID808 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID809 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID810 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID811 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID191_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [1:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid0 , nid1 , nid1 , nid1 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID812 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID813 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID192_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [5:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid0 , nid0 , nid0 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID814 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID815 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID816 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID817 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID818 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID819 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID193_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [5:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid0 , nid0 , nid0 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID820 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID821 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID822 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID823 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID824 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID825 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID194_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [0:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid0 , nid0 , nid0 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID826 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID195_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [2:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid0 , nid0 , nid0 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID827 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID828 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID829 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID196_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [4:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid0 , nid0 , nid0 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID830 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID831 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID832 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID833 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID834 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID197_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [2:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid0 , nid0 , nid0 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID835 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID836 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID837 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID198_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [2:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid0 , nid0 , nid0 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID838 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID839 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID840 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID199_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [6:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid0 , nid0 , nid0 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID841 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID842 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID843 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID844 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID845 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID846 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID847 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID200_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [0:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid0 , nid0 , nid1 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID848 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID201_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [1:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid0 , nid0 , nid1 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID849 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID850 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID202_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [4:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid0 , nid0 , nid1 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID851 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID852 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID853 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID854 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID855 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID203_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [2:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid0 , nid0 , nid1 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID856 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID857 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID858 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID204_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [5:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid0 , nid0 , nid1 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID859 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID860 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID861 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID862 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID863 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID864 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID205_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [2:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid0 , nid0 , nid1 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID865 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID866 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID867 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID206_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [2:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid0 , nid0 , nid1 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID868 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID869 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID870 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID207_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [1:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid0 , nid0 , nid1 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID871 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID872 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID208_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [4:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid0 , nid1 , nid0 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID873 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID874 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID875 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID876 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID877 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID209_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [1:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid0 , nid1 , nid0 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID878 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID879 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID210_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [5:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid0 , nid1 , nid0 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID880 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID881 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID882 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID883 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID884 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID885 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID211_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [5:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid0 , nid1 , nid0 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID886 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID887 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID888 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID889 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID890 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID891 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID212_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [1:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid0 , nid1 , nid0 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID892 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID893 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID213_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [1:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid0 , nid1 , nid0 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID894 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID895 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID214_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [6:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid0 , nid1 , nid0 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID896 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID897 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID898 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID899 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID900 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID901 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID902 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID215_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [0:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid0 , nid1 , nid0 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID903 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID216_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [5:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid0 , nid1 , nid1 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID904 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID905 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID906 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID907 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID908 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID909 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID217_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [3:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid0 , nid1 , nid1 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID910 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID911 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID912 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID913 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID218_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [1:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid0 , nid1 , nid1 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID914 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID915 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID219_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [2:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid0 , nid1 , nid1 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID916 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID917 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID918 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID220_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [4:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid0 , nid1 , nid1 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID919 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID920 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID921 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID922 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID923 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID221_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [2:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid0 , nid1 , nid1 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID924 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID925 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID926 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID222_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [0:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid0 , nid1 , nid1 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID927 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID223_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [2:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid0 , nid1 , nid1 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID928 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID929 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID930 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID224_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [6:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid1 , nid0 , nid0 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID931 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID932 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID933 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID934 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID935 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID936 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID937 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID225_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [4:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid1 , nid0 , nid0 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID938 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID939 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID940 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID941 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID942 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID226_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [4:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid1 , nid0 , nid0 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID943 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID944 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID945 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID946 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID947 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID227_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [0:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid1 , nid0 , nid0 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID948 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID228_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [1:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid1 , nid0 , nid0 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID949 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID950 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID229_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [5:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid1 , nid0 , nid0 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID951 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID952 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID953 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID954 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID955 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID956 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID230_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [2:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid1 , nid0 , nid0 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID957 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID958 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID959 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID231_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [2:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid1 , nid0 , nid0 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID960 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID961 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID962 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID232_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [0:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid1 , nid0 , nid1 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID963 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID233_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [5:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid1 , nid0 , nid1 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID964 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID965 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID966 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID967 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID968 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID969 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID234_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [0:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid1 , nid0 , nid1 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID970 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID235_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [2:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid1 , nid0 , nid1 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID971 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID972 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID973 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID236_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [1:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid1 , nid0 , nid1 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID974 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID975 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID237_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [3:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid1 , nid0 , nid1 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID976 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID977 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID978 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID979 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID238_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [6:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid1 , nid0 , nid1 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID980 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID981 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID982 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID983 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID984 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID985 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID986 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID239_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [4:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid1 , nid0 , nid1 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID987 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID988 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID989 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID990 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID991 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID240_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [0:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid1 , nid1 , nid0 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID992 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID241_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [3:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid1 , nid1 , nid0 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID993 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID994 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID995 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID996 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID242_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [3:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid1 , nid1 , nid0 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID997 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID998 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID999 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1000 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID243_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [2:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid1 , nid1 , nid0 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1001 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1002 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1003 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID244_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [3:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid1 , nid1 , nid0 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1004 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1005 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1006 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1007 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID245_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [2:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid1 , nid1 , nid0 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1008 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1009 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1010 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID246_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [4:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid1 , nid1 , nid0 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1011 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1012 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1013 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1014 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1015 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID247_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [4:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid1 , nid1 , nid0 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1016 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1017 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1018 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1019 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1020 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID248_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [1:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid1 , nid1 , nid1 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1021 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1022 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID249_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [6:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid1 , nid1 , nid1 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1023 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1024 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1025 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1026 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1027 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1028 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1029 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID250_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [0:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid1 , nid1 , nid1 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1030 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID251_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [4:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid1 , nid1 , nid1 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1031 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1032 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1033 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1034 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1035 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID252_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [0:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid1 , nid1 , nid1 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1036 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID253_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [1:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid1 , nid1 , nid1 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1037 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1038 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID254_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [4:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid1 , nid1 , nid1 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1039 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1040 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1041 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1042 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1043 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID255_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [0:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid0 , nid1 , nid1 , nid1 , nid1 , nid1 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1044 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID256_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [5:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid0 , nid0 , nid0 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1045 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1046 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1047 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1048 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1049 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1050 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID257_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [2:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid0 , nid0 , nid0 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1051 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1052 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1053 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID258_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [4:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid0 , nid0 , nid0 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1054 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1055 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1056 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1057 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1058 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID259_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [3:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid0 , nid0 , nid0 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1059 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1060 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1061 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1062 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID260_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [5:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid0 , nid0 , nid0 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1063 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1064 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1065 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1066 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1067 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1068 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID261_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [2:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid0 , nid0 , nid0 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1069 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1070 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1071 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID262_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [1:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid0 , nid0 , nid0 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1072 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1073 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID263_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [2:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid0 , nid0 , nid0 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1074 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1075 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1076 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID264_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [1:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid0 , nid0 , nid1 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1077 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1078 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID265_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [0:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid0 , nid0 , nid1 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1079 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID266_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [6:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid0 , nid0 , nid1 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1080 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1081 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1082 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1083 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1084 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1085 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1086 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID267_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [4:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid0 , nid0 , nid1 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1087 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1088 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1089 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1090 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1091 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID268_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [1:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid0 , nid0 , nid1 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1092 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1093 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID269_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [0:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid0 , nid0 , nid1 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1094 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID270_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [4:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid0 , nid0 , nid1 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1095 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1096 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1097 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1098 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1099 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID271_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [4:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid0 , nid0 , nid1 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1100 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1101 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1102 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1103 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1104 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID272_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [4:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid0 , nid1 , nid0 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1105 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1106 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1107 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1108 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1109 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID273_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [6:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid0 , nid1 , nid0 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1110 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1111 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1112 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1113 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1114 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1115 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1116 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID274_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [0:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid0 , nid1 , nid0 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1117 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID275_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [0:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid0 , nid1 , nid0 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1118 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID276_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [5:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid0 , nid1 , nid0 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1119 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1120 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1121 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1122 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1123 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1124 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID277_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [0:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid0 , nid1 , nid0 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1125 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID278_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [3:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid0 , nid1 , nid0 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1126 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1127 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1128 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1129 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID279_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [0:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid0 , nid1 , nid0 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1130 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID280_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [5:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid0 , nid1 , nid1 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1131 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1132 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1133 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1134 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1135 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1136 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID281_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [2:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid0 , nid1 , nid1 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1137 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1138 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1139 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID282_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [2:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid0 , nid1 , nid1 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1140 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1141 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1142 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID283_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [6:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid0 , nid1 , nid1 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1143 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1144 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1145 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1146 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1147 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1148 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1149 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID284_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [1:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid0 , nid1 , nid1 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1150 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1151 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID285_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [1:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid0 , nid1 , nid1 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1152 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1153 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID286_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [4:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid0 , nid1 , nid1 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1154 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1155 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1156 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1157 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1158 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID287_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [0:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid0 , nid1 , nid1 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1159 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID288_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [2:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid1 , nid0 , nid0 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1160 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1161 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1162 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID289_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [1:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid1 , nid0 , nid0 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1163 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1164 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID290_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [0:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid1 , nid0 , nid0 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1165 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID291_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [2:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid1 , nid0 , nid0 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1166 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1167 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1168 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID292_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [2:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid1 , nid0 , nid0 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1169 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1170 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1171 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID293_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [0:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid1 , nid0 , nid0 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1172 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID294_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [5:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid1 , nid0 , nid0 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1173 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1174 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1175 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1176 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1177 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1178 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID295_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [4:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid1 , nid0 , nid0 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1179 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1180 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1181 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1182 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1183 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID296_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [0:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid1 , nid0 , nid1 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1184 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID297_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [4:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid1 , nid0 , nid1 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1185 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1186 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1187 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1188 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1189 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID298_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [6:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid1 , nid0 , nid1 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1190 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1191 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1192 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1193 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1194 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1195 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1196 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID299_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [6:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid1 , nid0 , nid1 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1197 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1198 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1199 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1200 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1201 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1202 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1203 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID300_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [2:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid1 , nid0 , nid1 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1204 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1205 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1206 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID301_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [1:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid1 , nid0 , nid1 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1207 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1208 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID302_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [1:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid1 , nid0 , nid1 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1209 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1210 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID303_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [6:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid1 , nid0 , nid1 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1211 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1212 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1213 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1214 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1215 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1216 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1217 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID304_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [4:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid1 , nid1 , nid0 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1218 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1219 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1220 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1221 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1222 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID305_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [2:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid1 , nid1 , nid0 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1223 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1224 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1225 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID306_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [1:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid1 , nid1 , nid0 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1226 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1227 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID307_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [1:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid1 , nid1 , nid0 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1228 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1229 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID308_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [3:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid1 , nid1 , nid0 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1230 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1231 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1232 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1233 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID309_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [4:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid1 , nid1 , nid0 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1234 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1235 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1236 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1237 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1238 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID310_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [4:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid1 , nid1 , nid0 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1239 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1240 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1241 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1242 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1243 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID311_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [3:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid1 , nid1 , nid0 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1244 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1245 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1246 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1247 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID312_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [4:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid1 , nid1 , nid1 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1248 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1249 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1250 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1251 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1252 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID313_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [1:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid1 , nid1 , nid1 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1253 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1254 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID314_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [0:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid1 , nid1 , nid1 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1255 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID315_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [5:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid1 , nid1 , nid1 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1256 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1257 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1258 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1259 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1260 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1261 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID316_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [4:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid1 , nid1 , nid1 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1262 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1263 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1264 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1265 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1266 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID317_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [3:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid1 , nid1 , nid1 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1267 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1268 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1269 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1270 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID318_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [2:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid1 , nid1 , nid1 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1271 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1272 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1273 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID319_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [0:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid0 , nid1 , nid1 , nid1 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1274 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID320_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [6:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid0 , nid0 , nid0 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1275 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1276 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1277 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1278 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1279 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1280 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1281 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID321_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [0:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid0 , nid0 , nid0 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1282 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID322_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [6:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid0 , nid0 , nid0 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1283 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1284 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1285 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1286 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1287 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1288 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1289 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID323_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [2:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid0 , nid0 , nid0 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1290 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1291 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1292 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID324_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [6:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid0 , nid0 , nid0 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1293 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1294 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1295 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1296 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1297 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1298 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1299 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID325_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [1:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid0 , nid0 , nid0 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1300 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1301 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID326_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [4:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid0 , nid0 , nid0 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1302 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1303 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1304 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1305 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1306 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID327_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [2:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid0 , nid0 , nid0 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1307 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1308 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1309 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID328_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [5:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid0 , nid0 , nid1 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1310 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1311 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1312 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1313 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1314 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1315 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID329_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [6:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid0 , nid0 , nid1 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1316 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1317 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1318 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1319 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1320 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1321 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1322 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID330_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [4:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid0 , nid0 , nid1 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1323 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1324 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1325 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1326 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1327 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID331_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [5:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid0 , nid0 , nid1 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1328 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1329 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1330 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1331 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1332 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1333 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID332_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [5:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid0 , nid0 , nid1 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1334 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1335 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1336 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1337 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1338 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1339 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID333_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [3:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid0 , nid0 , nid1 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1340 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1341 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1342 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1343 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID334_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [2:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid0 , nid0 , nid1 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1344 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1345 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1346 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID335_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [4:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid0 , nid0 , nid1 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1347 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1348 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1349 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1350 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1351 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID336_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [3:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid0 , nid1 , nid0 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1352 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1353 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1354 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1355 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID337_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [2:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid0 , nid1 , nid0 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1356 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1357 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1358 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID338_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [0:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid0 , nid1 , nid0 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1359 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID339_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [2:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid0 , nid1 , nid0 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1360 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1361 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1362 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID340_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [4:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid0 , nid1 , nid0 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1363 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1364 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1365 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1366 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1367 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID341_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [5:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid0 , nid1 , nid0 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1368 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1369 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1370 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1371 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1372 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1373 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID342_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [2:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid0 , nid1 , nid0 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1374 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1375 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1376 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID343_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [0:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid0 , nid1 , nid0 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1377 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID344_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [3:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid0 , nid1 , nid1 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1378 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1379 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1380 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1381 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID345_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [4:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid0 , nid1 , nid1 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1382 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1383 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1384 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1385 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1386 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID346_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [6:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid0 , nid1 , nid1 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1387 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1388 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1389 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1390 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1391 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1392 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1393 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID347_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [2:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid0 , nid1 , nid1 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1394 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1395 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1396 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID348_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [1:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid0 , nid1 , nid1 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1397 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1398 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID349_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [1:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid0 , nid1 , nid1 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1399 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1400 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID350_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [5:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid0 , nid1 , nid1 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1401 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1402 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1403 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1404 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1405 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1406 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID351_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [1:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid0 , nid1 , nid1 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1407 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1408 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID352_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [0:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid1 , nid0 , nid0 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1409 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID353_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [3:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid1 , nid0 , nid0 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1410 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1411 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1412 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1413 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID354_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [6:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid1 , nid0 , nid0 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1414 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1415 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1416 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1417 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1418 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1419 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1420 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID355_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [3:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid1 , nid0 , nid0 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1421 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1422 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1423 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1424 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID356_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [4:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid1 , nid0 , nid0 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1425 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1426 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1427 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1428 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1429 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID357_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [0:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid1 , nid0 , nid0 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1430 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID358_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [3:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid1 , nid0 , nid0 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1431 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1432 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1433 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1434 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID359_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [5:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid1 , nid0 , nid0 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1435 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1436 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1437 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1438 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1439 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1440 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID360_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [5:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid1 , nid0 , nid1 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1441 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1442 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1443 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1444 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1445 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1446 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID361_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [4:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid1 , nid0 , nid1 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1447 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1448 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1449 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1450 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1451 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID362_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [2:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid1 , nid0 , nid1 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1452 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1453 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1454 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID363_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [2:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid1 , nid0 , nid1 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1455 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1456 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1457 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID364_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [4:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid1 , nid0 , nid1 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1458 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1459 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1460 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1461 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1462 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID365_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [2:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid1 , nid0 , nid1 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1463 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1464 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1465 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID366_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [0:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid1 , nid0 , nid1 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1466 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID367_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [5:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid1 , nid0 , nid1 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1467 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1468 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1469 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1470 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1471 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1472 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID368_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [5:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid1 , nid1 , nid0 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1473 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1474 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1475 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1476 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1477 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1478 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID369_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [4:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid1 , nid1 , nid0 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1479 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1480 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1481 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1482 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1483 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID370_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [4:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid1 , nid1 , nid0 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1484 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1485 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1486 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1487 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1488 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID371_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [6:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid1 , nid1 , nid0 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1489 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1490 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1491 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1492 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1493 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1494 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1495 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID372_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [3:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid1 , nid1 , nid0 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1496 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1497 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1498 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1499 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID373_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [1:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid1 , nid1 , nid0 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1500 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1501 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID374_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [5:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid1 , nid1 , nid0 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1502 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1503 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1504 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1505 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1506 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1507 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID375_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [1:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid1 , nid1 , nid0 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1508 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1509 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID376_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [3:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid1 , nid1 , nid1 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1510 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1511 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1512 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1513 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID377_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [3:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid1 , nid1 , nid1 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1514 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1515 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1516 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1517 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID378_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [4:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid1 , nid1 , nid1 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1518 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1519 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1520 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1521 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1522 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID379_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [3:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid1 , nid1 , nid1 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1523 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1524 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1525 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1526 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID380_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [1:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid1 , nid1 , nid1 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1527 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1528 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID381_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [4:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid1 , nid1 , nid1 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1529 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1530 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1531 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1532 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1533 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID382_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [2:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid1 , nid1 , nid1 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1534 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1535 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1536 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID383_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [2:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid1 , nid0 , nid1 , nid1 , nid1 , nid1 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1537 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1538 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1539 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID384_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [0:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid0 , nid0 , nid0 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1540 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID385_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [2:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid0 , nid0 , nid0 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1541 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1542 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1543 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID386_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [5:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid0 , nid0 , nid0 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1544 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1545 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1546 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1547 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1548 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1549 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID387_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [6:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid0 , nid0 , nid0 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1550 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1551 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1552 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1553 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1554 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1555 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1556 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID388_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [6:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid0 , nid0 , nid0 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1557 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1558 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1559 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1560 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1561 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1562 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1563 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID389_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [3:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid0 , nid0 , nid0 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1564 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1565 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1566 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1567 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID390_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [4:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid0 , nid0 , nid0 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1568 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1569 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1570 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1571 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1572 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID391_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [5:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid0 , nid0 , nid0 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1573 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1574 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1575 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1576 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1577 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1578 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID392_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [4:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid0 , nid0 , nid1 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1579 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1580 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1581 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1582 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1583 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID393_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [5:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid0 , nid0 , nid1 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1584 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1585 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1586 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1587 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1588 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1589 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID394_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [0:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid0 , nid0 , nid1 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1590 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID395_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [0:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid0 , nid0 , nid1 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1591 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID396_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [6:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid0 , nid0 , nid1 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1592 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1593 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1594 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1595 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1596 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1597 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1598 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID397_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [5:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid0 , nid0 , nid1 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1599 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1600 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1601 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1602 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1603 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1604 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID398_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [3:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid0 , nid0 , nid1 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1605 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1606 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1607 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1608 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID399_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [4:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid0 , nid0 , nid1 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1609 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1610 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1611 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1612 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1613 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID400_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [6:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid0 , nid1 , nid0 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1614 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1615 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1616 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1617 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1618 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1619 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1620 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID401_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [6:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid0 , nid1 , nid0 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1621 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1622 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1623 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1624 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1625 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1626 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1627 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID402_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [6:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid0 , nid1 , nid0 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1628 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1629 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1630 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1631 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1632 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1633 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1634 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID403_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [6:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid0 , nid1 , nid0 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1635 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1636 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1637 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1638 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1639 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1640 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1641 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID404_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [1:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid0 , nid1 , nid0 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1642 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1643 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID405_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [5:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid0 , nid1 , nid0 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1644 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1645 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1646 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1647 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1648 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1649 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID406_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [0:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid0 , nid1 , nid0 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1650 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID407_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [1:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid0 , nid1 , nid0 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1651 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1652 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID408_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [5:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid0 , nid1 , nid1 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1653 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1654 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1655 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1656 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1657 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1658 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID409_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [3:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid0 , nid1 , nid1 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1659 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1660 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1661 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1662 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID410_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [1:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid0 , nid1 , nid1 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1663 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1664 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID411_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [0:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid0 , nid1 , nid1 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1665 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID412_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [3:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid0 , nid1 , nid1 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1666 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1667 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1668 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1669 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID413_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [3:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid0 , nid1 , nid1 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1670 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1671 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1672 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1673 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID414_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [6:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid0 , nid1 , nid1 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1674 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1675 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1676 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1677 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1678 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1679 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1680 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID415_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [3:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid0 , nid1 , nid1 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1681 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1682 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1683 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1684 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID416_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [4:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid1 , nid0 , nid0 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1685 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1686 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1687 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1688 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1689 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID417_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [2:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid1 , nid0 , nid0 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1690 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1691 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1692 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID418_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [2:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid1 , nid0 , nid0 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1693 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1694 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1695 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID419_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [5:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid1 , nid0 , nid0 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1696 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1697 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1698 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1699 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1700 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1701 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID420_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [1:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid1 , nid0 , nid0 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1702 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1703 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID421_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [5:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid1 , nid0 , nid0 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1704 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1705 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1706 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1707 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1708 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1709 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID422_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [2:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid1 , nid0 , nid0 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1710 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1711 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1712 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID423_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [0:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid1 , nid0 , nid0 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1713 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID424_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [5:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid1 , nid0 , nid1 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1714 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1715 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1716 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1717 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1718 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1719 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID425_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [1:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid1 , nid0 , nid1 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1720 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1721 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID426_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [6:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid1 , nid0 , nid1 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1722 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1723 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1724 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1725 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1726 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1727 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1728 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID427_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [0:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid1 , nid0 , nid1 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1729 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID428_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [1:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid1 , nid0 , nid1 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1730 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1731 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID429_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [0:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid1 , nid0 , nid1 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1732 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID430_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [0:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid1 , nid0 , nid1 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1733 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID431_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [0:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid1 , nid0 , nid1 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1734 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID432_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [2:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid1 , nid1 , nid0 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1735 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1736 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1737 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID433_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [6:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid1 , nid1 , nid0 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1738 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1739 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1740 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1741 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1742 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1743 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1744 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID434_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [5:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid1 , nid1 , nid0 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1745 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1746 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1747 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1748 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1749 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1750 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID435_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [1:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid1 , nid1 , nid0 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1751 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1752 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID436_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [6:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid1 , nid1 , nid0 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1753 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1754 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1755 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1756 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1757 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1758 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1759 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID437_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [3:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid1 , nid1 , nid0 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1760 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1761 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1762 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1763 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID438_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [2:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid1 , nid1 , nid0 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1764 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1765 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1766 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID439_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [0:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid1 , nid1 , nid0 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1767 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID440_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [6:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid1 , nid1 , nid1 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1768 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1769 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1770 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1771 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1772 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1773 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1774 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID441_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [2:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid1 , nid1 , nid1 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1775 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1776 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1777 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID442_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [1:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid1 , nid1 , nid1 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1778 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1779 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID443_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [5:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid1 , nid1 , nid1 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1780 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1781 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1782 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1783 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1784 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1785 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID444_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [1:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid1 , nid1 , nid1 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1786 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1787 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID445_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [2:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid1 , nid1 , nid1 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1788 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1789 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1790 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID446_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [3:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid1 , nid1 , nid1 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1791 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1792 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1793 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1794 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID447_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [0:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid0 , nid1 , nid1 , nid1 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1795 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID448_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [2:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid0 , nid0 , nid0 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1796 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1797 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1798 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID449_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [6:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid0 , nid0 , nid0 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1799 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1800 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1801 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1802 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1803 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1804 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1805 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID450_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [3:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid0 , nid0 , nid0 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1806 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1807 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1808 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1809 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID451_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [0:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid0 , nid0 , nid0 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1810 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID452_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [1:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid0 , nid0 , nid0 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1811 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1812 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID453_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [4:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid0 , nid0 , nid0 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1813 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1814 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1815 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1816 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1817 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID454_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [4:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid0 , nid0 , nid0 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1818 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1819 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1820 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1821 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1822 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID455_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [6:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid0 , nid0 , nid0 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1823 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1824 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1825 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1826 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1827 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1828 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1829 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID456_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [1:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid0 , nid0 , nid1 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1830 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1831 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID457_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [5:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid0 , nid0 , nid1 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1832 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1833 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1834 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1835 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1836 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1837 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID458_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [6:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid0 , nid0 , nid1 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1838 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1839 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1840 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1841 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1842 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1843 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1844 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID459_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [4:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid0 , nid0 , nid1 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1845 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1846 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1847 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1848 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1849 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID460_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [6:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid0 , nid0 , nid1 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1850 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1851 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1852 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1853 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1854 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1855 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1856 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID461_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [0:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid0 , nid0 , nid1 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1857 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID462_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [5:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid0 , nid0 , nid1 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1858 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1859 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1860 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1861 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1862 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1863 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID463_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [0:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid0 , nid0 , nid1 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1864 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID464_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [3:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid0 , nid1 , nid0 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1865 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1866 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1867 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1868 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID465_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [6:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid0 , nid1 , nid0 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1869 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1870 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1871 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1872 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1873 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1874 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1875 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID466_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [3:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid0 , nid1 , nid0 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1876 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1877 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1878 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1879 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID467_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [4:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid0 , nid1 , nid0 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1880 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1881 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1882 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1883 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1884 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID468_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [0:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid0 , nid1 , nid0 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1885 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID469_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [3:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid0 , nid1 , nid0 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1886 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1887 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1888 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1889 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID470_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [1:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid0 , nid1 , nid0 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1890 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1891 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID471_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [3:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid0 , nid1 , nid0 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1892 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1893 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1894 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1895 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID472_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [5:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid0 , nid1 , nid1 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1896 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1897 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1898 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1899 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1900 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1901 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID473_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [1:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid0 , nid1 , nid1 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1902 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1903 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID474_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [1:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid0 , nid1 , nid1 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1904 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1905 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID475_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [6:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid0 , nid1 , nid1 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1906 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1907 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1908 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1909 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1910 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1911 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1912 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID476_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [4:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid0 , nid1 , nid1 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1913 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1914 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1915 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1916 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1917 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID477_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [0:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid0 , nid1 , nid1 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1918 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID478_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [6:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid0 , nid1 , nid1 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1919 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1920 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1921 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1922 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1923 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1924 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1925 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID479_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [3:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid0 , nid1 , nid1 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1926 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1927 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1928 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1929 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID480_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [4:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid1 , nid0 , nid0 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1930 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1931 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1932 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1933 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1934 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID481_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [1:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid1 , nid0 , nid0 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1935 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1936 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID482_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [2:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid1 , nid0 , nid0 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1937 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1938 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1939 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID483_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [2:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid1 , nid0 , nid0 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1940 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1941 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1942 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID484_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [1:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid1 , nid0 , nid0 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1943 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1944 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID485_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [0:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid1 , nid0 , nid0 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1945 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID486_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [0:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid1 , nid0 , nid0 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1946 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID487_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [0:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid1 , nid0 , nid0 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1947 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID488_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [6:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid1 , nid0 , nid1 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1948 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1949 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1950 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1951 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1952 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1953 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1954 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID489_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [1:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid1 , nid0 , nid1 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1955 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1956 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID490_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [3:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid1 , nid0 , nid1 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1957 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1958 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1959 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1960 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID491_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [2:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid1 , nid0 , nid1 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1961 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1962 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1963 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID492_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [4:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid1 , nid0 , nid1 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1964 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1965 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1966 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1967 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1968 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID493_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [6:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid1 , nid0 , nid1 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1969 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1970 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1971 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1972 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1973 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1974 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1975 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID494_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [2:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid1 , nid0 , nid1 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1976 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1977 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1978 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID495_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [2:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid1 , nid0 , nid1 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1979 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1980 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1981 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID496_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [3:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid1 , nid1 , nid0 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1982 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1983 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1984 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1985 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID497_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [5:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid1 , nid1 , nid0 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1986 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1987 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1988 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1989 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1990 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1991 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID498_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [4:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid1 , nid1 , nid0 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1992 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1993 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1994 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1995 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1996 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID499_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [3:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid1 , nid1 , nid0 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID1997 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1998 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID1999 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID2000 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID500_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [0:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid1 , nid1 , nid0 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID2001 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID501_INDEGREE4 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [3:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE4_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid1 , nid1 , nid0 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID2002 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID2003 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID2004 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID2005 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID502_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [5:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid1 , nid1 , nid0 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID2006 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID2007 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID2008 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID2009 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID2010 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID2011 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID503_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [6:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid1 , nid1 , nid0 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID2012 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID2013 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID2014 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID2015 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID2016 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID2017 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID2018 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID504_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [0:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid1 , nid1 , nid1 , nid0 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID2019 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID505_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [6:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid1 , nid1 , nid1 , nid0 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID2020 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID2021 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID2022 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID2023 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID2024 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID2025 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID2026 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID506_INDEGREE6 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [5:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE6_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid1 , nid1 , nid1 , nid0 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID2027 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID2028 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID2029 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID2030 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID2031 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID2032 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID507_INDEGREE5 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [4:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE5_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid1 , nid1 , nid1 , nid0 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID2033 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID2034 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID2035 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID2036 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID2037 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID508_INDEGREE7 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [6:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE7_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid1 , nid1 , nid1 , nid1 , nid0 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID2038 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID2039 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID2040 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID2041 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID2042 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID2043 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID2044 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID509_INDEGREE1 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [0:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE1_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid1 , nid1 , nid1 , nid1 , nid0 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID2045 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID510_INDEGREE3 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [2:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE3_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid1 , nid1 , nid1 , nid1 , nid1 , nid0  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID2046 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID2047 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid0 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID2048 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module Node_NID511_INDEGREE2 ( InEdges, OutEdge, PathAddr, PathData, Start, Clk );
input  [1:0] InEdges;
output [0:0] OutEdge;
input  [8:0] PathAddr;
output [2:0] PathData;
input Start, Clk;

    wire nid0, nid1;
    NodeAux_INDEGREE2_SOURCE0 nodeAux ( .Nid({nid1 , nid1 , nid1 , nid1 , nid1 , nid1 , nid1 , nid1 , nid1  }),
        .InEdges(InEdges), .OutEdge(OutEdge),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(nid1 ) );
    VMW_PULLDOWN U4 ( .Z(nid0 ) );
endmodule

module Edge_EID2049 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule

module Edge_EID2050 (InEdge, OutEdge, WeightAddr, WeightData, Clk );
input  [0:0] InEdge;
input  [11:0] WeightAddr;
output [0:0] OutEdge;
input  [0:0] WeightData;
input  Clk;
    wire eid0, eid1;
    EdgeAux edgeAux ( .Eid({eid1 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid0 , eid1 , eid0  }),
        .InEdge(InEdge), .OutEdge(OutEdge),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    VMW_PULLUP U3 ( .Z(eid1 ) );
    VMW_PULLDOWN U4 ( .Z(eid0 ) );
endmodule


module graph ( WeightAddr, WeightData, PathAddr, PathData, Start, Clk );
input  [11:0] WeightAddr;
input  [0:0] WeightData;
input  [8:0] PathAddr;
output [2:0] PathData;
input  Start, Clk;
    wire [0:0] In0;
    wire [0:0] Out0;
    wire [5:0] In1;
    wire [0:0] Out1;
    wire [3:0] In2;
    wire [0:0] Out2;
    wire [5:0] In3;
    wire [0:0] Out3;
    wire [6:0] In4;
    wire [0:0] Out4;
    wire [0:0] In5;
    wire [0:0] Out5;
    wire [6:0] In6;
    wire [0:0] Out6;
    wire [3:0] In7;
    wire [0:0] Out7;
    wire [6:0] In8;
    wire [0:0] Out8;
    wire [5:0] In9;
    wire [0:0] Out9;
    wire [5:0] In10;
    wire [0:0] Out10;
    wire [3:0] In11;
    wire [0:0] Out11;
    wire [5:0] In12;
    wire [0:0] Out12;
    wire [5:0] In13;
    wire [0:0] Out13;
    wire [4:0] In14;
    wire [0:0] Out14;
    wire [1:0] In15;
    wire [0:0] Out15;
    wire [3:0] In16;
    wire [0:0] Out16;
    wire [1:0] In17;
    wire [0:0] Out17;
    wire [5:0] In18;
    wire [0:0] Out18;
    wire [6:0] In19;
    wire [0:0] Out19;
    wire [6:0] In20;
    wire [0:0] Out20;
    wire [3:0] In21;
    wire [0:0] Out21;
    wire [6:0] In22;
    wire [0:0] Out22;
    wire [3:0] In23;
    wire [0:0] Out23;
    wire [0:0] In24;
    wire [0:0] Out24;
    wire [6:0] In25;
    wire [0:0] Out25;
    wire [4:0] In26;
    wire [0:0] Out26;
    wire [5:0] In27;
    wire [0:0] Out27;
    wire [0:0] In28;
    wire [0:0] Out28;
    wire [2:0] In29;
    wire [0:0] Out29;
    wire [0:0] In30;
    wire [0:0] Out30;
    wire [5:0] In31;
    wire [0:0] Out31;
    wire [1:0] In32;
    wire [0:0] Out32;
    wire [6:0] In33;
    wire [0:0] Out33;
    wire [2:0] In34;
    wire [0:0] Out34;
    wire [5:0] In35;
    wire [0:0] Out35;
    wire [4:0] In36;
    wire [0:0] Out36;
    wire [6:0] In37;
    wire [0:0] Out37;
    wire [5:0] In38;
    wire [0:0] Out38;
    wire [1:0] In39;
    wire [0:0] Out39;
    wire [4:0] In40;
    wire [0:0] Out40;
    wire [0:0] In41;
    wire [0:0] Out41;
    wire [4:0] In42;
    wire [0:0] Out42;
    wire [2:0] In43;
    wire [0:0] Out43;
    wire [0:0] In44;
    wire [0:0] Out44;
    wire [2:0] In45;
    wire [0:0] Out45;
    wire [2:0] In46;
    wire [0:0] Out46;
    wire [3:0] In47;
    wire [0:0] Out47;
    wire [0:0] In48;
    wire [0:0] Out48;
    wire [6:0] In49;
    wire [0:0] Out49;
    wire [4:0] In50;
    wire [0:0] Out50;
    wire [6:0] In51;
    wire [0:0] Out51;
    wire [3:0] In52;
    wire [0:0] Out52;
    wire [0:0] In53;
    wire [0:0] Out53;
    wire [0:0] In54;
    wire [0:0] Out54;
    wire [4:0] In55;
    wire [0:0] Out55;
    wire [4:0] In56;
    wire [0:0] Out56;
    wire [2:0] In57;
    wire [0:0] Out57;
    wire [5:0] In58;
    wire [0:0] Out58;
    wire [2:0] In59;
    wire [0:0] Out59;
    wire [2:0] In60;
    wire [0:0] Out60;
    wire [0:0] In61;
    wire [0:0] Out61;
    wire [4:0] In62;
    wire [0:0] Out62;
    wire [4:0] In63;
    wire [0:0] Out63;
    wire [1:0] In64;
    wire [0:0] Out64;
    wire [4:0] In65;
    wire [0:0] Out65;
    wire [4:0] In66;
    wire [0:0] Out66;
    wire [1:0] In67;
    wire [0:0] Out67;
    wire [4:0] In68;
    wire [0:0] Out68;
    wire [3:0] In69;
    wire [0:0] Out69;
    wire [0:0] In70;
    wire [0:0] Out70;
    wire [3:0] In71;
    wire [0:0] Out71;
    wire [6:0] In72;
    wire [0:0] Out72;
    wire [0:0] In73;
    wire [0:0] Out73;
    wire [4:0] In74;
    wire [0:0] Out74;
    wire [1:0] In75;
    wire [0:0] Out75;
    wire [2:0] In76;
    wire [0:0] Out76;
    wire [4:0] In77;
    wire [0:0] Out77;
    wire [6:0] In78;
    wire [0:0] Out78;
    wire [2:0] In79;
    wire [0:0] Out79;
    wire [6:0] In80;
    wire [0:0] Out80;
    wire [0:0] In81;
    wire [0:0] Out81;
    wire [0:0] In82;
    wire [0:0] Out82;
    wire [5:0] In83;
    wire [0:0] Out83;
    wire [4:0] In84;
    wire [0:0] Out84;
    wire [1:0] In85;
    wire [0:0] Out85;
    wire [0:0] In86;
    wire [0:0] Out86;
    wire [2:0] In87;
    wire [0:0] Out87;
    wire [4:0] In88;
    wire [0:0] Out88;
    wire [6:0] In89;
    wire [0:0] Out89;
    wire [2:0] In90;
    wire [0:0] Out90;
    wire [5:0] In91;
    wire [0:0] Out91;
    wire [5:0] In92;
    wire [0:0] Out92;
    wire [2:0] In93;
    wire [0:0] Out93;
    wire [0:0] In94;
    wire [0:0] Out94;
    wire [5:0] In95;
    wire [0:0] Out95;
    wire [4:0] In96;
    wire [0:0] Out96;
    wire [3:0] In97;
    wire [0:0] Out97;
    wire [5:0] In98;
    wire [0:0] Out98;
    wire [4:0] In99;
    wire [0:0] Out99;
    wire [3:0] In100;
    wire [0:0] Out100;
    wire [3:0] In101;
    wire [0:0] Out101;
    wire [3:0] In102;
    wire [0:0] Out102;
    wire [2:0] In103;
    wire [0:0] Out103;
    wire [4:0] In104;
    wire [0:0] Out104;
    wire [2:0] In105;
    wire [0:0] Out105;
    wire [6:0] In106;
    wire [0:0] Out106;
    wire [4:0] In107;
    wire [0:0] Out107;
    wire [4:0] In108;
    wire [0:0] Out108;
    wire [1:0] In109;
    wire [0:0] Out109;
    wire [4:0] In110;
    wire [0:0] Out110;
    wire [6:0] In111;
    wire [0:0] Out111;
    wire [4:0] In112;
    wire [0:0] Out112;
    wire [1:0] In113;
    wire [0:0] Out113;
    wire [2:0] In114;
    wire [0:0] Out114;
    wire [3:0] In115;
    wire [0:0] Out115;
    wire [6:0] In116;
    wire [0:0] Out116;
    wire [1:0] In117;
    wire [0:0] Out117;
    wire [1:0] In118;
    wire [0:0] Out118;
    wire [6:0] In119;
    wire [0:0] Out119;
    wire [5:0] In120;
    wire [0:0] Out120;
    wire [5:0] In121;
    wire [0:0] Out121;
    wire [6:0] In122;
    wire [0:0] Out122;
    wire [0:0] In123;
    wire [0:0] Out123;
    wire [2:0] In124;
    wire [0:0] Out124;
    wire [0:0] In125;
    wire [0:0] Out125;
    wire [4:0] In126;
    wire [0:0] Out126;
    wire [5:0] In127;
    wire [0:0] Out127;
    wire [2:0] In128;
    wire [0:0] Out128;
    wire [2:0] In129;
    wire [0:0] Out129;
    wire [1:0] In130;
    wire [0:0] Out130;
    wire [3:0] In131;
    wire [0:0] Out131;
    wire [4:0] In132;
    wire [0:0] Out132;
    wire [6:0] In133;
    wire [0:0] Out133;
    wire [2:0] In134;
    wire [0:0] Out134;
    wire [6:0] In135;
    wire [0:0] Out135;
    wire [4:0] In136;
    wire [0:0] Out136;
    wire [2:0] In137;
    wire [0:0] Out137;
    wire [0:0] In138;
    wire [0:0] Out138;
    wire [1:0] In139;
    wire [0:0] Out139;
    wire [3:0] In140;
    wire [0:0] Out140;
    wire [6:0] In141;
    wire [0:0] Out141;
    wire [0:0] In142;
    wire [0:0] Out142;
    wire [5:0] In143;
    wire [0:0] Out143;
    wire [5:0] In144;
    wire [0:0] Out144;
    wire [2:0] In145;
    wire [0:0] Out145;
    wire [2:0] In146;
    wire [0:0] Out146;
    wire [4:0] In147;
    wire [0:0] Out147;
    wire [6:0] In148;
    wire [0:0] Out148;
    wire [3:0] In149;
    wire [0:0] Out149;
    wire [5:0] In150;
    wire [0:0] Out150;
    wire [2:0] In151;
    wire [0:0] Out151;
    wire [6:0] In152;
    wire [0:0] Out152;
    wire [3:0] In153;
    wire [0:0] Out153;
    wire [6:0] In154;
    wire [0:0] Out154;
    wire [0:0] In155;
    wire [0:0] Out155;
    wire [4:0] In156;
    wire [0:0] Out156;
    wire [6:0] In157;
    wire [0:0] Out157;
    wire [1:0] In158;
    wire [0:0] Out158;
    wire [6:0] In159;
    wire [0:0] Out159;
    wire [6:0] In160;
    wire [0:0] Out160;
    wire [3:0] In161;
    wire [0:0] Out161;
    wire [1:0] In162;
    wire [0:0] Out162;
    wire [6:0] In163;
    wire [0:0] Out163;
    wire [4:0] In164;
    wire [0:0] Out164;
    wire [0:0] In165;
    wire [0:0] Out165;
    wire [0:0] In166;
    wire [0:0] Out166;
    wire [5:0] In167;
    wire [0:0] Out167;
    wire [0:0] In168;
    wire [0:0] Out168;
    wire [3:0] In169;
    wire [0:0] Out169;
    wire [4:0] In170;
    wire [0:0] Out170;
    wire [4:0] In171;
    wire [0:0] Out171;
    wire [6:0] In172;
    wire [0:0] Out172;
    wire [1:0] In173;
    wire [0:0] Out173;
    wire [1:0] In174;
    wire [0:0] Out174;
    wire [0:0] In175;
    wire [0:0] Out175;
    wire [4:0] In176;
    wire [0:0] Out176;
    wire [0:0] In177;
    wire [0:0] Out177;
    wire [4:0] In178;
    wire [0:0] Out178;
    wire [6:0] In179;
    wire [0:0] Out179;
    wire [5:0] In180;
    wire [0:0] Out180;
    wire [6:0] In181;
    wire [0:0] Out181;
    wire [6:0] In182;
    wire [0:0] Out182;
    wire [3:0] In183;
    wire [0:0] Out183;
    wire [6:0] In184;
    wire [0:0] Out184;
    wire [0:0] In185;
    wire [0:0] Out185;
    wire [0:0] In186;
    wire [0:0] Out186;
    wire [2:0] In187;
    wire [0:0] Out187;
    wire [4:0] In188;
    wire [0:0] Out188;
    wire [6:0] In189;
    wire [0:0] Out189;
    wire [6:0] In190;
    wire [0:0] Out190;
    wire [1:0] In191;
    wire [0:0] Out191;
    wire [5:0] In192;
    wire [0:0] Out192;
    wire [5:0] In193;
    wire [0:0] Out193;
    wire [0:0] In194;
    wire [0:0] Out194;
    wire [2:0] In195;
    wire [0:0] Out195;
    wire [4:0] In196;
    wire [0:0] Out196;
    wire [2:0] In197;
    wire [0:0] Out197;
    wire [2:0] In198;
    wire [0:0] Out198;
    wire [6:0] In199;
    wire [0:0] Out199;
    wire [0:0] In200;
    wire [0:0] Out200;
    wire [1:0] In201;
    wire [0:0] Out201;
    wire [4:0] In202;
    wire [0:0] Out202;
    wire [2:0] In203;
    wire [0:0] Out203;
    wire [5:0] In204;
    wire [0:0] Out204;
    wire [2:0] In205;
    wire [0:0] Out205;
    wire [2:0] In206;
    wire [0:0] Out206;
    wire [1:0] In207;
    wire [0:0] Out207;
    wire [4:0] In208;
    wire [0:0] Out208;
    wire [1:0] In209;
    wire [0:0] Out209;
    wire [5:0] In210;
    wire [0:0] Out210;
    wire [5:0] In211;
    wire [0:0] Out211;
    wire [1:0] In212;
    wire [0:0] Out212;
    wire [1:0] In213;
    wire [0:0] Out213;
    wire [6:0] In214;
    wire [0:0] Out214;
    wire [0:0] In215;
    wire [0:0] Out215;
    wire [5:0] In216;
    wire [0:0] Out216;
    wire [3:0] In217;
    wire [0:0] Out217;
    wire [1:0] In218;
    wire [0:0] Out218;
    wire [2:0] In219;
    wire [0:0] Out219;
    wire [4:0] In220;
    wire [0:0] Out220;
    wire [2:0] In221;
    wire [0:0] Out221;
    wire [0:0] In222;
    wire [0:0] Out222;
    wire [2:0] In223;
    wire [0:0] Out223;
    wire [6:0] In224;
    wire [0:0] Out224;
    wire [4:0] In225;
    wire [0:0] Out225;
    wire [4:0] In226;
    wire [0:0] Out226;
    wire [0:0] In227;
    wire [0:0] Out227;
    wire [1:0] In228;
    wire [0:0] Out228;
    wire [5:0] In229;
    wire [0:0] Out229;
    wire [2:0] In230;
    wire [0:0] Out230;
    wire [2:0] In231;
    wire [0:0] Out231;
    wire [0:0] In232;
    wire [0:0] Out232;
    wire [5:0] In233;
    wire [0:0] Out233;
    wire [0:0] In234;
    wire [0:0] Out234;
    wire [2:0] In235;
    wire [0:0] Out235;
    wire [1:0] In236;
    wire [0:0] Out236;
    wire [3:0] In237;
    wire [0:0] Out237;
    wire [6:0] In238;
    wire [0:0] Out238;
    wire [4:0] In239;
    wire [0:0] Out239;
    wire [0:0] In240;
    wire [0:0] Out240;
    wire [3:0] In241;
    wire [0:0] Out241;
    wire [3:0] In242;
    wire [0:0] Out242;
    wire [2:0] In243;
    wire [0:0] Out243;
    wire [3:0] In244;
    wire [0:0] Out244;
    wire [2:0] In245;
    wire [0:0] Out245;
    wire [4:0] In246;
    wire [0:0] Out246;
    wire [4:0] In247;
    wire [0:0] Out247;
    wire [1:0] In248;
    wire [0:0] Out248;
    wire [6:0] In249;
    wire [0:0] Out249;
    wire [0:0] In250;
    wire [0:0] Out250;
    wire [4:0] In251;
    wire [0:0] Out251;
    wire [0:0] In252;
    wire [0:0] Out252;
    wire [1:0] In253;
    wire [0:0] Out253;
    wire [4:0] In254;
    wire [0:0] Out254;
    wire [0:0] In255;
    wire [0:0] Out255;
    wire [5:0] In256;
    wire [0:0] Out256;
    wire [2:0] In257;
    wire [0:0] Out257;
    wire [4:0] In258;
    wire [0:0] Out258;
    wire [3:0] In259;
    wire [0:0] Out259;
    wire [5:0] In260;
    wire [0:0] Out260;
    wire [2:0] In261;
    wire [0:0] Out261;
    wire [1:0] In262;
    wire [0:0] Out262;
    wire [2:0] In263;
    wire [0:0] Out263;
    wire [1:0] In264;
    wire [0:0] Out264;
    wire [0:0] In265;
    wire [0:0] Out265;
    wire [6:0] In266;
    wire [0:0] Out266;
    wire [4:0] In267;
    wire [0:0] Out267;
    wire [1:0] In268;
    wire [0:0] Out268;
    wire [0:0] In269;
    wire [0:0] Out269;
    wire [4:0] In270;
    wire [0:0] Out270;
    wire [4:0] In271;
    wire [0:0] Out271;
    wire [4:0] In272;
    wire [0:0] Out272;
    wire [6:0] In273;
    wire [0:0] Out273;
    wire [0:0] In274;
    wire [0:0] Out274;
    wire [0:0] In275;
    wire [0:0] Out275;
    wire [5:0] In276;
    wire [0:0] Out276;
    wire [0:0] In277;
    wire [0:0] Out277;
    wire [3:0] In278;
    wire [0:0] Out278;
    wire [0:0] In279;
    wire [0:0] Out279;
    wire [5:0] In280;
    wire [0:0] Out280;
    wire [2:0] In281;
    wire [0:0] Out281;
    wire [2:0] In282;
    wire [0:0] Out282;
    wire [6:0] In283;
    wire [0:0] Out283;
    wire [1:0] In284;
    wire [0:0] Out284;
    wire [1:0] In285;
    wire [0:0] Out285;
    wire [4:0] In286;
    wire [0:0] Out286;
    wire [0:0] In287;
    wire [0:0] Out287;
    wire [2:0] In288;
    wire [0:0] Out288;
    wire [1:0] In289;
    wire [0:0] Out289;
    wire [0:0] In290;
    wire [0:0] Out290;
    wire [2:0] In291;
    wire [0:0] Out291;
    wire [2:0] In292;
    wire [0:0] Out292;
    wire [0:0] In293;
    wire [0:0] Out293;
    wire [5:0] In294;
    wire [0:0] Out294;
    wire [4:0] In295;
    wire [0:0] Out295;
    wire [0:0] In296;
    wire [0:0] Out296;
    wire [4:0] In297;
    wire [0:0] Out297;
    wire [6:0] In298;
    wire [0:0] Out298;
    wire [6:0] In299;
    wire [0:0] Out299;
    wire [2:0] In300;
    wire [0:0] Out300;
    wire [1:0] In301;
    wire [0:0] Out301;
    wire [1:0] In302;
    wire [0:0] Out302;
    wire [6:0] In303;
    wire [0:0] Out303;
    wire [4:0] In304;
    wire [0:0] Out304;
    wire [2:0] In305;
    wire [0:0] Out305;
    wire [1:0] In306;
    wire [0:0] Out306;
    wire [1:0] In307;
    wire [0:0] Out307;
    wire [3:0] In308;
    wire [0:0] Out308;
    wire [4:0] In309;
    wire [0:0] Out309;
    wire [4:0] In310;
    wire [0:0] Out310;
    wire [3:0] In311;
    wire [0:0] Out311;
    wire [4:0] In312;
    wire [0:0] Out312;
    wire [1:0] In313;
    wire [0:0] Out313;
    wire [0:0] In314;
    wire [0:0] Out314;
    wire [5:0] In315;
    wire [0:0] Out315;
    wire [4:0] In316;
    wire [0:0] Out316;
    wire [3:0] In317;
    wire [0:0] Out317;
    wire [2:0] In318;
    wire [0:0] Out318;
    wire [0:0] In319;
    wire [0:0] Out319;
    wire [6:0] In320;
    wire [0:0] Out320;
    wire [0:0] In321;
    wire [0:0] Out321;
    wire [6:0] In322;
    wire [0:0] Out322;
    wire [2:0] In323;
    wire [0:0] Out323;
    wire [6:0] In324;
    wire [0:0] Out324;
    wire [1:0] In325;
    wire [0:0] Out325;
    wire [4:0] In326;
    wire [0:0] Out326;
    wire [2:0] In327;
    wire [0:0] Out327;
    wire [5:0] In328;
    wire [0:0] Out328;
    wire [6:0] In329;
    wire [0:0] Out329;
    wire [4:0] In330;
    wire [0:0] Out330;
    wire [5:0] In331;
    wire [0:0] Out331;
    wire [5:0] In332;
    wire [0:0] Out332;
    wire [3:0] In333;
    wire [0:0] Out333;
    wire [2:0] In334;
    wire [0:0] Out334;
    wire [4:0] In335;
    wire [0:0] Out335;
    wire [3:0] In336;
    wire [0:0] Out336;
    wire [2:0] In337;
    wire [0:0] Out337;
    wire [0:0] In338;
    wire [0:0] Out338;
    wire [2:0] In339;
    wire [0:0] Out339;
    wire [4:0] In340;
    wire [0:0] Out340;
    wire [5:0] In341;
    wire [0:0] Out341;
    wire [2:0] In342;
    wire [0:0] Out342;
    wire [0:0] In343;
    wire [0:0] Out343;
    wire [3:0] In344;
    wire [0:0] Out344;
    wire [4:0] In345;
    wire [0:0] Out345;
    wire [6:0] In346;
    wire [0:0] Out346;
    wire [2:0] In347;
    wire [0:0] Out347;
    wire [1:0] In348;
    wire [0:0] Out348;
    wire [1:0] In349;
    wire [0:0] Out349;
    wire [5:0] In350;
    wire [0:0] Out350;
    wire [1:0] In351;
    wire [0:0] Out351;
    wire [0:0] In352;
    wire [0:0] Out352;
    wire [3:0] In353;
    wire [0:0] Out353;
    wire [6:0] In354;
    wire [0:0] Out354;
    wire [3:0] In355;
    wire [0:0] Out355;
    wire [4:0] In356;
    wire [0:0] Out356;
    wire [0:0] In357;
    wire [0:0] Out357;
    wire [3:0] In358;
    wire [0:0] Out358;
    wire [5:0] In359;
    wire [0:0] Out359;
    wire [5:0] In360;
    wire [0:0] Out360;
    wire [4:0] In361;
    wire [0:0] Out361;
    wire [2:0] In362;
    wire [0:0] Out362;
    wire [2:0] In363;
    wire [0:0] Out363;
    wire [4:0] In364;
    wire [0:0] Out364;
    wire [2:0] In365;
    wire [0:0] Out365;
    wire [0:0] In366;
    wire [0:0] Out366;
    wire [5:0] In367;
    wire [0:0] Out367;
    wire [5:0] In368;
    wire [0:0] Out368;
    wire [4:0] In369;
    wire [0:0] Out369;
    wire [4:0] In370;
    wire [0:0] Out370;
    wire [6:0] In371;
    wire [0:0] Out371;
    wire [3:0] In372;
    wire [0:0] Out372;
    wire [1:0] In373;
    wire [0:0] Out373;
    wire [5:0] In374;
    wire [0:0] Out374;
    wire [1:0] In375;
    wire [0:0] Out375;
    wire [3:0] In376;
    wire [0:0] Out376;
    wire [3:0] In377;
    wire [0:0] Out377;
    wire [4:0] In378;
    wire [0:0] Out378;
    wire [3:0] In379;
    wire [0:0] Out379;
    wire [1:0] In380;
    wire [0:0] Out380;
    wire [4:0] In381;
    wire [0:0] Out381;
    wire [2:0] In382;
    wire [0:0] Out382;
    wire [2:0] In383;
    wire [0:0] Out383;
    wire [0:0] In384;
    wire [0:0] Out384;
    wire [2:0] In385;
    wire [0:0] Out385;
    wire [5:0] In386;
    wire [0:0] Out386;
    wire [6:0] In387;
    wire [0:0] Out387;
    wire [6:0] In388;
    wire [0:0] Out388;
    wire [3:0] In389;
    wire [0:0] Out389;
    wire [4:0] In390;
    wire [0:0] Out390;
    wire [5:0] In391;
    wire [0:0] Out391;
    wire [4:0] In392;
    wire [0:0] Out392;
    wire [5:0] In393;
    wire [0:0] Out393;
    wire [0:0] In394;
    wire [0:0] Out394;
    wire [0:0] In395;
    wire [0:0] Out395;
    wire [6:0] In396;
    wire [0:0] Out396;
    wire [5:0] In397;
    wire [0:0] Out397;
    wire [3:0] In398;
    wire [0:0] Out398;
    wire [4:0] In399;
    wire [0:0] Out399;
    wire [6:0] In400;
    wire [0:0] Out400;
    wire [6:0] In401;
    wire [0:0] Out401;
    wire [6:0] In402;
    wire [0:0] Out402;
    wire [6:0] In403;
    wire [0:0] Out403;
    wire [1:0] In404;
    wire [0:0] Out404;
    wire [5:0] In405;
    wire [0:0] Out405;
    wire [0:0] In406;
    wire [0:0] Out406;
    wire [1:0] In407;
    wire [0:0] Out407;
    wire [5:0] In408;
    wire [0:0] Out408;
    wire [3:0] In409;
    wire [0:0] Out409;
    wire [1:0] In410;
    wire [0:0] Out410;
    wire [0:0] In411;
    wire [0:0] Out411;
    wire [3:0] In412;
    wire [0:0] Out412;
    wire [3:0] In413;
    wire [0:0] Out413;
    wire [6:0] In414;
    wire [0:0] Out414;
    wire [3:0] In415;
    wire [0:0] Out415;
    wire [4:0] In416;
    wire [0:0] Out416;
    wire [2:0] In417;
    wire [0:0] Out417;
    wire [2:0] In418;
    wire [0:0] Out418;
    wire [5:0] In419;
    wire [0:0] Out419;
    wire [1:0] In420;
    wire [0:0] Out420;
    wire [5:0] In421;
    wire [0:0] Out421;
    wire [2:0] In422;
    wire [0:0] Out422;
    wire [0:0] In423;
    wire [0:0] Out423;
    wire [5:0] In424;
    wire [0:0] Out424;
    wire [1:0] In425;
    wire [0:0] Out425;
    wire [6:0] In426;
    wire [0:0] Out426;
    wire [0:0] In427;
    wire [0:0] Out427;
    wire [1:0] In428;
    wire [0:0] Out428;
    wire [0:0] In429;
    wire [0:0] Out429;
    wire [0:0] In430;
    wire [0:0] Out430;
    wire [0:0] In431;
    wire [0:0] Out431;
    wire [2:0] In432;
    wire [0:0] Out432;
    wire [6:0] In433;
    wire [0:0] Out433;
    wire [5:0] In434;
    wire [0:0] Out434;
    wire [1:0] In435;
    wire [0:0] Out435;
    wire [6:0] In436;
    wire [0:0] Out436;
    wire [3:0] In437;
    wire [0:0] Out437;
    wire [2:0] In438;
    wire [0:0] Out438;
    wire [0:0] In439;
    wire [0:0] Out439;
    wire [6:0] In440;
    wire [0:0] Out440;
    wire [2:0] In441;
    wire [0:0] Out441;
    wire [1:0] In442;
    wire [0:0] Out442;
    wire [5:0] In443;
    wire [0:0] Out443;
    wire [1:0] In444;
    wire [0:0] Out444;
    wire [2:0] In445;
    wire [0:0] Out445;
    wire [3:0] In446;
    wire [0:0] Out446;
    wire [0:0] In447;
    wire [0:0] Out447;
    wire [2:0] In448;
    wire [0:0] Out448;
    wire [6:0] In449;
    wire [0:0] Out449;
    wire [3:0] In450;
    wire [0:0] Out450;
    wire [0:0] In451;
    wire [0:0] Out451;
    wire [1:0] In452;
    wire [0:0] Out452;
    wire [4:0] In453;
    wire [0:0] Out453;
    wire [4:0] In454;
    wire [0:0] Out454;
    wire [6:0] In455;
    wire [0:0] Out455;
    wire [1:0] In456;
    wire [0:0] Out456;
    wire [5:0] In457;
    wire [0:0] Out457;
    wire [6:0] In458;
    wire [0:0] Out458;
    wire [4:0] In459;
    wire [0:0] Out459;
    wire [6:0] In460;
    wire [0:0] Out460;
    wire [0:0] In461;
    wire [0:0] Out461;
    wire [5:0] In462;
    wire [0:0] Out462;
    wire [0:0] In463;
    wire [0:0] Out463;
    wire [3:0] In464;
    wire [0:0] Out464;
    wire [6:0] In465;
    wire [0:0] Out465;
    wire [3:0] In466;
    wire [0:0] Out466;
    wire [4:0] In467;
    wire [0:0] Out467;
    wire [0:0] In468;
    wire [0:0] Out468;
    wire [3:0] In469;
    wire [0:0] Out469;
    wire [1:0] In470;
    wire [0:0] Out470;
    wire [3:0] In471;
    wire [0:0] Out471;
    wire [5:0] In472;
    wire [0:0] Out472;
    wire [1:0] In473;
    wire [0:0] Out473;
    wire [1:0] In474;
    wire [0:0] Out474;
    wire [6:0] In475;
    wire [0:0] Out475;
    wire [4:0] In476;
    wire [0:0] Out476;
    wire [0:0] In477;
    wire [0:0] Out477;
    wire [6:0] In478;
    wire [0:0] Out478;
    wire [3:0] In479;
    wire [0:0] Out479;
    wire [4:0] In480;
    wire [0:0] Out480;
    wire [1:0] In481;
    wire [0:0] Out481;
    wire [2:0] In482;
    wire [0:0] Out482;
    wire [2:0] In483;
    wire [0:0] Out483;
    wire [1:0] In484;
    wire [0:0] Out484;
    wire [0:0] In485;
    wire [0:0] Out485;
    wire [0:0] In486;
    wire [0:0] Out486;
    wire [0:0] In487;
    wire [0:0] Out487;
    wire [6:0] In488;
    wire [0:0] Out488;
    wire [1:0] In489;
    wire [0:0] Out489;
    wire [3:0] In490;
    wire [0:0] Out490;
    wire [2:0] In491;
    wire [0:0] Out491;
    wire [4:0] In492;
    wire [0:0] Out492;
    wire [6:0] In493;
    wire [0:0] Out493;
    wire [2:0] In494;
    wire [0:0] Out494;
    wire [2:0] In495;
    wire [0:0] Out495;
    wire [3:0] In496;
    wire [0:0] Out496;
    wire [5:0] In497;
    wire [0:0] Out497;
    wire [4:0] In498;
    wire [0:0] Out498;
    wire [3:0] In499;
    wire [0:0] Out499;
    wire [0:0] In500;
    wire [0:0] Out500;
    wire [3:0] In501;
    wire [0:0] Out501;
    wire [5:0] In502;
    wire [0:0] Out502;
    wire [6:0] In503;
    wire [0:0] Out503;
    wire [0:0] In504;
    wire [0:0] Out504;
    wire [6:0] In505;
    wire [0:0] Out505;
    wire [5:0] In506;
    wire [0:0] Out506;
    wire [4:0] In507;
    wire [0:0] Out507;
    wire [6:0] In508;
    wire [0:0] Out508;
    wire [0:0] In509;
    wire [0:0] Out509;
    wire [2:0] In510;
    wire [0:0] Out510;
    wire [1:0] In511;
    wire [0:0] Out511;

    Node_NID0_INDEGREE1 n0 ( .InEdges(In0), .OutEdge(Out0),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID0 e0 ( .InEdge(Out435), .OutEdge(In0[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID1_INDEGREE6 n1 ( .InEdges(In1), .OutEdge(Out1),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1 e1 ( .InEdge(Out143), .OutEdge(In1[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID2 e2 ( .InEdge(Out452), .OutEdge(In1[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID3 e3 ( .InEdge(Out171), .OutEdge(In1[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID4 e4 ( .InEdge(Out155), .OutEdge(In1[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID5 e5 ( .InEdge(Out509), .OutEdge(In1[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID6 e6 ( .InEdge(Out400), .OutEdge(In1[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID2_INDEGREE4 n2 ( .InEdges(In2), .OutEdge(Out2),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID7 e7 ( .InEdge(Out177), .OutEdge(In2[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID8 e8 ( .InEdge(Out91), .OutEdge(In2[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID9 e9 ( .InEdge(Out94), .OutEdge(In2[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID10 e10 ( .InEdge(Out304), .OutEdge(In2[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID3_INDEGREE6 n3 ( .InEdges(In3), .OutEdge(Out3),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID11 e11 ( .InEdge(Out27), .OutEdge(In3[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID12 e12 ( .InEdge(Out130), .OutEdge(In3[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID13 e13 ( .InEdge(Out102), .OutEdge(In3[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID14 e14 ( .InEdge(Out293), .OutEdge(In3[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID15 e15 ( .InEdge(Out15), .OutEdge(In3[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID16 e16 ( .InEdge(Out429), .OutEdge(In3[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID4_INDEGREE7 n4 ( .InEdges(In4), .OutEdge(Out4),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID17 e17 ( .InEdge(Out368), .OutEdge(In4[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID18 e18 ( .InEdge(Out258), .OutEdge(In4[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID19 e19 ( .InEdge(Out106), .OutEdge(In4[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID20 e20 ( .InEdge(Out25), .OutEdge(In4[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID21 e21 ( .InEdge(Out475), .OutEdge(In4[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID22 e22 ( .InEdge(Out419), .OutEdge(In4[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID23 e23 ( .InEdge(Out190), .OutEdge(In4[6:6]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID5_INDEGREE1 n5 ( .InEdges(In5), .OutEdge(Out5),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID24 e24 ( .InEdge(Out312), .OutEdge(In5[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID6_INDEGREE7 n6 ( .InEdges(In6), .OutEdge(Out6),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID25 e25 ( .InEdge(Out458), .OutEdge(In6[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID26 e26 ( .InEdge(Out42), .OutEdge(In6[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID27 e27 ( .InEdge(Out352), .OutEdge(In6[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID28 e28 ( .InEdge(Out394), .OutEdge(In6[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID29 e29 ( .InEdge(Out144), .OutEdge(In6[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID30 e30 ( .InEdge(Out405), .OutEdge(In6[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID31 e31 ( .InEdge(Out206), .OutEdge(In6[6:6]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID7_INDEGREE4 n7 ( .InEdges(In7), .OutEdge(Out7),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID32 e32 ( .InEdge(Out423), .OutEdge(In7[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID33 e33 ( .InEdge(Out323), .OutEdge(In7[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID34 e34 ( .InEdge(Out495), .OutEdge(In7[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID35 e35 ( .InEdge(Out115), .OutEdge(In7[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID8_INDEGREE7 n8 ( .InEdges(In8), .OutEdge(Out8),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID36 e36 ( .InEdge(Out349), .OutEdge(In8[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID37 e37 ( .InEdge(Out453), .OutEdge(In8[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID38 e38 ( .InEdge(Out390), .OutEdge(In8[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID39 e39 ( .InEdge(Out501), .OutEdge(In8[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID40 e40 ( .InEdge(Out457), .OutEdge(In8[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID41 e41 ( .InEdge(Out487), .OutEdge(In8[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID42 e42 ( .InEdge(Out331), .OutEdge(In8[6:6]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID9_INDEGREE6 n9 ( .InEdges(In9), .OutEdge(Out9),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID43 e43 ( .InEdge(Out109), .OutEdge(In9[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID44 e44 ( .InEdge(Out51), .OutEdge(In9[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID45 e45 ( .InEdge(Out322), .OutEdge(In9[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID46 e46 ( .InEdge(Out510), .OutEdge(In9[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID47 e47 ( .InEdge(Out219), .OutEdge(In9[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID48 e48 ( .InEdge(Out12), .OutEdge(In9[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID10_INDEGREE6 n10 ( .InEdges(In10), .OutEdge(Out10),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID49 e49 ( .InEdge(Out170), .OutEdge(In10[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID50 e50 ( .InEdge(Out88), .OutEdge(In10[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID51 e51 ( .InEdge(Out30), .OutEdge(In10[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID52 e52 ( .InEdge(Out117), .OutEdge(In10[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID53 e53 ( .InEdge(Out287), .OutEdge(In10[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID54 e54 ( .InEdge(Out367), .OutEdge(In10[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID11_INDEGREE4 n11 ( .InEdges(In11), .OutEdge(Out11),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID55 e55 ( .InEdge(Out493), .OutEdge(In11[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID56 e56 ( .InEdge(Out444), .OutEdge(In11[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID57 e57 ( .InEdge(Out403), .OutEdge(In11[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID58 e58 ( .InEdge(Out342), .OutEdge(In11[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID12_INDEGREE6 n12 ( .InEdges(In12), .OutEdge(Out12),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID59 e59 ( .InEdge(Out194), .OutEdge(In12[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID60 e60 ( .InEdge(Out63), .OutEdge(In12[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID61 e61 ( .InEdge(Out379), .OutEdge(In12[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID62 e62 ( .InEdge(Out272), .OutEdge(In12[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID63 e63 ( .InEdge(Out442), .OutEdge(In12[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID64 e64 ( .InEdge(Out153), .OutEdge(In12[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID13_INDEGREE6 n13 ( .InEdges(In13), .OutEdge(Out13),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID65 e65 ( .InEdge(Out322), .OutEdge(In13[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID66 e66 ( .InEdge(Out188), .OutEdge(In13[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID67 e67 ( .InEdge(Out14), .OutEdge(In13[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID68 e68 ( .InEdge(Out104), .OutEdge(In13[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID69 e69 ( .InEdge(Out302), .OutEdge(In13[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID70 e70 ( .InEdge(Out240), .OutEdge(In13[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID14_INDEGREE5 n14 ( .InEdges(In14), .OutEdge(Out14),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID71 e71 ( .InEdge(Out392), .OutEdge(In14[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID72 e72 ( .InEdge(Out269), .OutEdge(In14[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID73 e73 ( .InEdge(Out196), .OutEdge(In14[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID74 e74 ( .InEdge(Out324), .OutEdge(In14[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID75 e75 ( .InEdge(Out285), .OutEdge(In14[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID15_INDEGREE2 n15 ( .InEdges(In15), .OutEdge(Out15),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID76 e76 ( .InEdge(Out230), .OutEdge(In15[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID77 e77 ( .InEdge(Out84), .OutEdge(In15[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID16_INDEGREE4 n16 ( .InEdges(In16), .OutEdge(Out16),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID78 e78 ( .InEdge(Out418), .OutEdge(In16[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID79 e79 ( .InEdge(Out166), .OutEdge(In16[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID80 e80 ( .InEdge(Out270), .OutEdge(In16[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID81 e81 ( .InEdge(Out460), .OutEdge(In16[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID17_INDEGREE2 n17 ( .InEdges(In17), .OutEdge(Out17),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID82 e82 ( .InEdge(Out497), .OutEdge(In17[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID83 e83 ( .InEdge(Out159), .OutEdge(In17[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID18_INDEGREE6 n18 ( .InEdges(In18), .OutEdge(Out18),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID84 e84 ( .InEdge(Out49), .OutEdge(In18[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID85 e85 ( .InEdge(Out471), .OutEdge(In18[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID86 e86 ( .InEdge(Out476), .OutEdge(In18[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID87 e87 ( .InEdge(Out407), .OutEdge(In18[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID88 e88 ( .InEdge(Out257), .OutEdge(In18[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID89 e89 ( .InEdge(Out361), .OutEdge(In18[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID19_INDEGREE7 n19 ( .InEdges(In19), .OutEdge(Out19),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID90 e90 ( .InEdge(Out381), .OutEdge(In19[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID91 e91 ( .InEdge(Out418), .OutEdge(In19[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID92 e92 ( .InEdge(Out419), .OutEdge(In19[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID93 e93 ( .InEdge(Out346), .OutEdge(In19[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID94 e94 ( .InEdge(Out447), .OutEdge(In19[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID95 e95 ( .InEdge(Out281), .OutEdge(In19[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID96 e96 ( .InEdge(Out325), .OutEdge(In19[6:6]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID20_INDEGREE7 n20 ( .InEdges(In20), .OutEdge(Out20),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID97 e97 ( .InEdge(Out219), .OutEdge(In20[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID98 e98 ( .InEdge(Out359), .OutEdge(In20[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID99 e99 ( .InEdge(Out254), .OutEdge(In20[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID100 e100 ( .InEdge(Out432), .OutEdge(In20[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID101 e101 ( .InEdge(Out281), .OutEdge(In20[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID102 e102 ( .InEdge(Out354), .OutEdge(In20[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID103 e103 ( .InEdge(Out67), .OutEdge(In20[6:6]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID21_INDEGREE4 n21 ( .InEdges(In21), .OutEdge(Out21),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID104 e104 ( .InEdge(Out226), .OutEdge(In21[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID105 e105 ( .InEdge(Out158), .OutEdge(In21[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID106 e106 ( .InEdge(Out54), .OutEdge(In21[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID107 e107 ( .InEdge(Out61), .OutEdge(In21[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID22_INDEGREE7 n22 ( .InEdges(In22), .OutEdge(Out22),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID108 e108 ( .InEdge(Out59), .OutEdge(In22[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID109 e109 ( .InEdge(Out300), .OutEdge(In22[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID110 e110 ( .InEdge(Out311), .OutEdge(In22[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID111 e111 ( .InEdge(Out392), .OutEdge(In22[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID112 e112 ( .InEdge(Out316), .OutEdge(In22[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID113 e113 ( .InEdge(Out485), .OutEdge(In22[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID114 e114 ( .InEdge(Out190), .OutEdge(In22[6:6]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID23_INDEGREE4 n23 ( .InEdges(In23), .OutEdge(Out23),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID115 e115 ( .InEdge(Out434), .OutEdge(In23[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID116 e116 ( .InEdge(Out55), .OutEdge(In23[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID117 e117 ( .InEdge(Out230), .OutEdge(In23[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID118 e118 ( .InEdge(Out295), .OutEdge(In23[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID24_INDEGREE1 n24 ( .InEdges(In24), .OutEdge(Out24),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID119 e119 ( .InEdge(Out175), .OutEdge(In24[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID25_INDEGREE7 n25 ( .InEdges(In25), .OutEdge(Out25),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID120 e120 ( .InEdge(Out48), .OutEdge(In25[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID121 e121 ( .InEdge(Out412), .OutEdge(In25[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID122 e122 ( .InEdge(Out433), .OutEdge(In25[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID123 e123 ( .InEdge(Out121), .OutEdge(In25[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID124 e124 ( .InEdge(Out464), .OutEdge(In25[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID125 e125 ( .InEdge(Out107), .OutEdge(In25[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID126 e126 ( .InEdge(Out130), .OutEdge(In25[6:6]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID26_INDEGREE5 n26 ( .InEdges(In26), .OutEdge(Out26),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID127 e127 ( .InEdge(Out18), .OutEdge(In26[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID128 e128 ( .InEdge(Out38), .OutEdge(In26[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID129 e129 ( .InEdge(Out178), .OutEdge(In26[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID130 e130 ( .InEdge(Out443), .OutEdge(In26[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID131 e131 ( .InEdge(Out347), .OutEdge(In26[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID27_INDEGREE6 n27 ( .InEdges(In27), .OutEdge(Out27),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID132 e132 ( .InEdge(Out304), .OutEdge(In27[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID133 e133 ( .InEdge(Out109), .OutEdge(In27[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID134 e134 ( .InEdge(Out11), .OutEdge(In27[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID135 e135 ( .InEdge(Out227), .OutEdge(In27[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID136 e136 ( .InEdge(Out458), .OutEdge(In27[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID137 e137 ( .InEdge(Out30), .OutEdge(In27[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID28_INDEGREE1 n28 ( .InEdges(In28), .OutEdge(Out28),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID138 e138 ( .InEdge(Out346), .OutEdge(In28[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID29_INDEGREE3 n29 ( .InEdges(In29), .OutEdge(Out29),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID139 e139 ( .InEdge(Out52), .OutEdge(In29[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID140 e140 ( .InEdge(Out75), .OutEdge(In29[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID141 e141 ( .InEdge(Out439), .OutEdge(In29[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID30_INDEGREE1 n30 ( .InEdges(In30), .OutEdge(Out30),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID142 e142 ( .InEdge(Out414), .OutEdge(In30[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID31_INDEGREE6 n31 ( .InEdges(In31), .OutEdge(Out31),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID143 e143 ( .InEdge(Out218), .OutEdge(In31[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID144 e144 ( .InEdge(Out63), .OutEdge(In31[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID145 e145 ( .InEdge(Out274), .OutEdge(In31[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID146 e146 ( .InEdge(Out464), .OutEdge(In31[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID147 e147 ( .InEdge(Out443), .OutEdge(In31[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID148 e148 ( .InEdge(Out135), .OutEdge(In31[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID32_INDEGREE2 n32 ( .InEdges(In32), .OutEdge(Out32),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID149 e149 ( .InEdge(Out460), .OutEdge(In32[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID150 e150 ( .InEdge(Out112), .OutEdge(In32[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID33_INDEGREE7 n33 ( .InEdges(In33), .OutEdge(Out33),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID151 e151 ( .InEdge(Out5), .OutEdge(In33[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID152 e152 ( .InEdge(Out402), .OutEdge(In33[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID153 e153 ( .InEdge(Out445), .OutEdge(In33[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID154 e154 ( .InEdge(Out45), .OutEdge(In33[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID155 e155 ( .InEdge(Out485), .OutEdge(In33[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID156 e156 ( .InEdge(Out229), .OutEdge(In33[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID157 e157 ( .InEdge(Out246), .OutEdge(In33[6:6]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID34_INDEGREE3 n34 ( .InEdges(In34), .OutEdge(Out34),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID158 e158 ( .InEdge(Out131), .OutEdge(In34[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID159 e159 ( .InEdge(Out411), .OutEdge(In34[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID160 e160 ( .InEdge(Out101), .OutEdge(In34[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID35_INDEGREE6 n35 ( .InEdges(In35), .OutEdge(Out35),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID161 e161 ( .InEdge(Out254), .OutEdge(In35[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID162 e162 ( .InEdge(Out271), .OutEdge(In35[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID163 e163 ( .InEdge(Out427), .OutEdge(In35[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID164 e164 ( .InEdge(Out367), .OutEdge(In35[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID165 e165 ( .InEdge(Out423), .OutEdge(In35[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID166 e166 ( .InEdge(Out236), .OutEdge(In35[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID36_INDEGREE5 n36 ( .InEdges(In36), .OutEdge(Out36),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID167 e167 ( .InEdge(Out226), .OutEdge(In36[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID168 e168 ( .InEdge(Out475), .OutEdge(In36[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID169 e169 ( .InEdge(Out225), .OutEdge(In36[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID170 e170 ( .InEdge(Out189), .OutEdge(In36[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID171 e171 ( .InEdge(Out308), .OutEdge(In36[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID37_INDEGREE7 n37 ( .InEdges(In37), .OutEdge(Out37),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID172 e172 ( .InEdge(Out143), .OutEdge(In37[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID173 e173 ( .InEdge(Out125), .OutEdge(In37[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID174 e174 ( .InEdge(Out488), .OutEdge(In37[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID175 e175 ( .InEdge(Out341), .OutEdge(In37[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID176 e176 ( .InEdge(Out273), .OutEdge(In37[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID177 e177 ( .InEdge(Out214), .OutEdge(In37[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID178 e178 ( .InEdge(Out254), .OutEdge(In37[6:6]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID38_INDEGREE6 n38 ( .InEdges(In38), .OutEdge(Out38),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID179 e179 ( .InEdge(Out356), .OutEdge(In38[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID180 e180 ( .InEdge(Out337), .OutEdge(In38[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID181 e181 ( .InEdge(Out47), .OutEdge(In38[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID182 e182 ( .InEdge(Out205), .OutEdge(In38[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID183 e183 ( .InEdge(Out19), .OutEdge(In38[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID184 e184 ( .InEdge(Out282), .OutEdge(In38[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID39_INDEGREE2 n39 ( .InEdges(In39), .OutEdge(Out39),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID185 e185 ( .InEdge(Out54), .OutEdge(In39[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID186 e186 ( .InEdge(Out477), .OutEdge(In39[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID40_INDEGREE5 n40 ( .InEdges(In40), .OutEdge(Out40),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID187 e187 ( .InEdge(Out300), .OutEdge(In40[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID188 e188 ( .InEdge(Out16), .OutEdge(In40[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID189 e189 ( .InEdge(Out480), .OutEdge(In40[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID190 e190 ( .InEdge(Out168), .OutEdge(In40[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID191 e191 ( .InEdge(Out113), .OutEdge(In40[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID41_INDEGREE1 n41 ( .InEdges(In41), .OutEdge(Out41),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID192 e192 ( .InEdge(Out175), .OutEdge(In41[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID42_INDEGREE5 n42 ( .InEdges(In42), .OutEdge(Out42),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID193 e193 ( .InEdge(Out57), .OutEdge(In42[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID194 e194 ( .InEdge(Out176), .OutEdge(In42[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID195 e195 ( .InEdge(Out131), .OutEdge(In42[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID196 e196 ( .InEdge(Out261), .OutEdge(In42[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID197 e197 ( .InEdge(Out266), .OutEdge(In42[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID43_INDEGREE3 n43 ( .InEdges(In43), .OutEdge(Out43),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID198 e198 ( .InEdge(Out438), .OutEdge(In43[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID199 e199 ( .InEdge(Out156), .OutEdge(In43[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID200 e200 ( .InEdge(Out363), .OutEdge(In43[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID44_INDEGREE1 n44 ( .InEdges(In44), .OutEdge(Out44),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID201 e201 ( .InEdge(Out213), .OutEdge(In44[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID45_INDEGREE3 n45 ( .InEdges(In45), .OutEdge(Out45),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID202 e202 ( .InEdge(Out268), .OutEdge(In45[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID203 e203 ( .InEdge(Out59), .OutEdge(In45[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID204 e204 ( .InEdge(Out35), .OutEdge(In45[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID46_INDEGREE3 n46 ( .InEdges(In46), .OutEdge(Out46),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID205 e205 ( .InEdge(Out63), .OutEdge(In46[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID206 e206 ( .InEdge(Out476), .OutEdge(In46[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID207 e207 ( .InEdge(Out23), .OutEdge(In46[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID47_INDEGREE4 n47 ( .InEdges(In47), .OutEdge(Out47),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID208 e208 ( .InEdge(Out36), .OutEdge(In47[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID209 e209 ( .InEdge(Out251), .OutEdge(In47[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID210 e210 ( .InEdge(Out18), .OutEdge(In47[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID211 e211 ( .InEdge(Out311), .OutEdge(In47[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID48_INDEGREE1 n48 ( .InEdges(In48), .OutEdge(Out48),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID212 e212 ( .InEdge(Out10), .OutEdge(In48[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID49_INDEGREE7 n49 ( .InEdges(In49), .OutEdge(Out49),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID213 e213 ( .InEdge(Out433), .OutEdge(In49[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID214 e214 ( .InEdge(Out169), .OutEdge(In49[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID215 e215 ( .InEdge(Out264), .OutEdge(In49[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID216 e216 ( .InEdge(Out283), .OutEdge(In49[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID217 e217 ( .InEdge(Out258), .OutEdge(In49[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID218 e218 ( .InEdge(Out381), .OutEdge(In49[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID219 e219 ( .InEdge(Out15), .OutEdge(In49[6:6]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID50_INDEGREE5 n50 ( .InEdges(In50), .OutEdge(Out50),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID220 e220 ( .InEdge(Out190), .OutEdge(In50[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID221 e221 ( .InEdge(Out272), .OutEdge(In50[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID222 e222 ( .InEdge(Out235), .OutEdge(In50[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID223 e223 ( .InEdge(Out118), .OutEdge(In50[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID224 e224 ( .InEdge(Out358), .OutEdge(In50[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID51_INDEGREE7 n51 ( .InEdges(In51), .OutEdge(Out51),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID225 e225 ( .InEdge(Out382), .OutEdge(In51[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID226 e226 ( .InEdge(Out437), .OutEdge(In51[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID227 e227 ( .InEdge(Out159), .OutEdge(In51[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID228 e228 ( .InEdge(Out54), .OutEdge(In51[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID229 e229 ( .InEdge(Out460), .OutEdge(In51[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID230 e230 ( .InEdge(Out288), .OutEdge(In51[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID231 e231 ( .InEdge(Out347), .OutEdge(In51[6:6]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID52_INDEGREE4 n52 ( .InEdges(In52), .OutEdge(Out52),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID232 e232 ( .InEdge(Out338), .OutEdge(In52[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID233 e233 ( .InEdge(Out359), .OutEdge(In52[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID234 e234 ( .InEdge(Out56), .OutEdge(In52[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID235 e235 ( .InEdge(Out215), .OutEdge(In52[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID53_INDEGREE1 n53 ( .InEdges(In53), .OutEdge(Out53),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID236 e236 ( .InEdge(Out382), .OutEdge(In53[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID54_INDEGREE1 n54 ( .InEdges(In54), .OutEdge(Out54),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID237 e237 ( .InEdge(Out17), .OutEdge(In54[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID55_INDEGREE5 n55 ( .InEdges(In55), .OutEdge(Out55),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID238 e238 ( .InEdge(Out18), .OutEdge(In55[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID239 e239 ( .InEdge(Out271), .OutEdge(In55[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID240 e240 ( .InEdge(Out459), .OutEdge(In55[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID241 e241 ( .InEdge(Out419), .OutEdge(In55[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID242 e242 ( .InEdge(Out252), .OutEdge(In55[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID56_INDEGREE5 n56 ( .InEdges(In56), .OutEdge(Out56),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID243 e243 ( .InEdge(Out308), .OutEdge(In56[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID244 e244 ( .InEdge(Out93), .OutEdge(In56[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID245 e245 ( .InEdge(Out123), .OutEdge(In56[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID246 e246 ( .InEdge(Out257), .OutEdge(In56[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID247 e247 ( .InEdge(Out305), .OutEdge(In56[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID57_INDEGREE3 n57 ( .InEdges(In57), .OutEdge(Out57),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID248 e248 ( .InEdge(Out102), .OutEdge(In57[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID249 e249 ( .InEdge(Out244), .OutEdge(In57[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID250 e250 ( .InEdge(Out112), .OutEdge(In57[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID58_INDEGREE6 n58 ( .InEdges(In58), .OutEdge(Out58),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID251 e251 ( .InEdge(Out330), .OutEdge(In58[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID252 e252 ( .InEdge(Out268), .OutEdge(In58[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID253 e253 ( .InEdge(Out109), .OutEdge(In58[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID254 e254 ( .InEdge(Out259), .OutEdge(In58[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID255 e255 ( .InEdge(Out403), .OutEdge(In58[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID256 e256 ( .InEdge(Out300), .OutEdge(In58[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID59_INDEGREE3 n59 ( .InEdges(In59), .OutEdge(Out59),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID257 e257 ( .InEdge(Out238), .OutEdge(In59[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID258 e258 ( .InEdge(Out152), .OutEdge(In59[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID259 e259 ( .InEdge(Out272), .OutEdge(In59[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID60_INDEGREE3 n60 ( .InEdges(In60), .OutEdge(Out60),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID260 e260 ( .InEdge(Out169), .OutEdge(In60[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID261 e261 ( .InEdge(Out41), .OutEdge(In60[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID262 e262 ( .InEdge(Out418), .OutEdge(In60[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID61_INDEGREE1 n61 ( .InEdges(In61), .OutEdge(Out61),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID263 e263 ( .InEdge(Out202), .OutEdge(In61[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID62_INDEGREE5 n62 ( .InEdges(In62), .OutEdge(Out62),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID264 e264 ( .InEdge(Out375), .OutEdge(In62[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID265 e265 ( .InEdge(Out422), .OutEdge(In62[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID266 e266 ( .InEdge(Out231), .OutEdge(In62[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID267 e267 ( .InEdge(Out54), .OutEdge(In62[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID268 e268 ( .InEdge(Out129), .OutEdge(In62[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID63_INDEGREE5 n63 ( .InEdges(In63), .OutEdge(Out63),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID269 e269 ( .InEdge(Out237), .OutEdge(In63[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID270 e270 ( .InEdge(Out432), .OutEdge(In63[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID271 e271 ( .InEdge(Out221), .OutEdge(In63[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID272 e272 ( .InEdge(Out74), .OutEdge(In63[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID273 e273 ( .InEdge(Out183), .OutEdge(In63[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID64_INDEGREE2 n64 ( .InEdges(In64), .OutEdge(Out64),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID274 e274 ( .InEdge(Out420), .OutEdge(In64[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID275 e275 ( .InEdge(Out28), .OutEdge(In64[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID65_INDEGREE5 n65 ( .InEdges(In65), .OutEdge(Out65),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID276 e276 ( .InEdge(Out80), .OutEdge(In65[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID277 e277 ( .InEdge(Out151), .OutEdge(In65[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID278 e278 ( .InEdge(Out271), .OutEdge(In65[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID279 e279 ( .InEdge(Out415), .OutEdge(In65[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID280 e280 ( .InEdge(Out174), .OutEdge(In65[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID66_INDEGREE5 n66 ( .InEdges(In66), .OutEdge(Out66),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID281 e281 ( .InEdge(Out131), .OutEdge(In66[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID282 e282 ( .InEdge(Out496), .OutEdge(In66[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID283 e283 ( .InEdge(Out399), .OutEdge(In66[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID284 e284 ( .InEdge(Out23), .OutEdge(In66[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID285 e285 ( .InEdge(Out272), .OutEdge(In66[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID67_INDEGREE2 n67 ( .InEdges(In67), .OutEdge(Out67),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID286 e286 ( .InEdge(Out445), .OutEdge(In67[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID287 e287 ( .InEdge(Out367), .OutEdge(In67[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID68_INDEGREE5 n68 ( .InEdges(In68), .OutEdge(Out68),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID288 e288 ( .InEdge(Out44), .OutEdge(In68[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID289 e289 ( .InEdge(Out378), .OutEdge(In68[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID290 e290 ( .InEdge(Out470), .OutEdge(In68[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID291 e291 ( .InEdge(Out58), .OutEdge(In68[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID292 e292 ( .InEdge(Out511), .OutEdge(In68[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID69_INDEGREE4 n69 ( .InEdges(In69), .OutEdge(Out69),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID293 e293 ( .InEdge(Out275), .OutEdge(In69[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID294 e294 ( .InEdge(Out236), .OutEdge(In69[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID295 e295 ( .InEdge(Out113), .OutEdge(In69[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID296 e296 ( .InEdge(Out239), .OutEdge(In69[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID70_INDEGREE1 n70 ( .InEdges(In70), .OutEdge(Out70),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID297 e297 ( .InEdge(Out50), .OutEdge(In70[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID71_INDEGREE4 n71 ( .InEdges(In71), .OutEdge(Out71),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID298 e298 ( .InEdge(Out159), .OutEdge(In71[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID299 e299 ( .InEdge(Out469), .OutEdge(In71[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID300 e300 ( .InEdge(Out280), .OutEdge(In71[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID301 e301 ( .InEdge(Out174), .OutEdge(In71[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID72_INDEGREE7 n72 ( .InEdges(In72), .OutEdge(Out72),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID302 e302 ( .InEdge(Out129), .OutEdge(In72[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID303 e303 ( .InEdge(Out102), .OutEdge(In72[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID304 e304 ( .InEdge(Out229), .OutEdge(In72[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID305 e305 ( .InEdge(Out169), .OutEdge(In72[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID306 e306 ( .InEdge(Out283), .OutEdge(In72[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID307 e307 ( .InEdge(Out400), .OutEdge(In72[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID308 e308 ( .InEdge(Out131), .OutEdge(In72[6:6]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID73_INDEGREE1 n73 ( .InEdges(In73), .OutEdge(Out73),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID309 e309 ( .InEdge(Out305), .OutEdge(In73[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID74_INDEGREE5 n74 ( .InEdges(In74), .OutEdge(Out74),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID310 e310 ( .InEdge(Out413), .OutEdge(In74[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID311 e311 ( .InEdge(Out292), .OutEdge(In74[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID312 e312 ( .InEdge(Out223), .OutEdge(In74[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID313 e313 ( .InEdge(Out113), .OutEdge(In74[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID314 e314 ( .InEdge(Out301), .OutEdge(In74[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID75_INDEGREE2 n75 ( .InEdges(In75), .OutEdge(Out75),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID315 e315 ( .InEdge(Out268), .OutEdge(In75[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID316 e316 ( .InEdge(Out182), .OutEdge(In75[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID76_INDEGREE3 n76 ( .InEdges(In76), .OutEdge(Out76),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID317 e317 ( .InEdge(Out495), .OutEdge(In76[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID318 e318 ( .InEdge(Out379), .OutEdge(In76[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID319 e319 ( .InEdge(Out180), .OutEdge(In76[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID77_INDEGREE5 n77 ( .InEdges(In77), .OutEdge(Out77),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID320 e320 ( .InEdge(Out19), .OutEdge(In77[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID321 e321 ( .InEdge(Out152), .OutEdge(In77[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID322 e322 ( .InEdge(Out190), .OutEdge(In77[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID323 e323 ( .InEdge(Out407), .OutEdge(In77[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID324 e324 ( .InEdge(Out273), .OutEdge(In77[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID78_INDEGREE7 n78 ( .InEdges(In78), .OutEdge(Out78),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID325 e325 ( .InEdge(Out340), .OutEdge(In78[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID326 e326 ( .InEdge(Out375), .OutEdge(In78[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID327 e327 ( .InEdge(Out177), .OutEdge(In78[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID328 e328 ( .InEdge(Out453), .OutEdge(In78[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID329 e329 ( .InEdge(Out66), .OutEdge(In78[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID330 e330 ( .InEdge(Out39), .OutEdge(In78[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID331 e331 ( .InEdge(Out194), .OutEdge(In78[6:6]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID79_INDEGREE3 n79 ( .InEdges(In79), .OutEdge(Out79),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID332 e332 ( .InEdge(Out422), .OutEdge(In79[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID333 e333 ( .InEdge(Out130), .OutEdge(In79[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID334 e334 ( .InEdge(Out296), .OutEdge(In79[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID80_INDEGREE7 n80 ( .InEdges(In80), .OutEdge(Out80),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID335 e335 ( .InEdge(Out389), .OutEdge(In80[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID336 e336 ( .InEdge(Out50), .OutEdge(In80[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID337 e337 ( .InEdge(Out222), .OutEdge(In80[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID338 e338 ( .InEdge(Out328), .OutEdge(In80[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID339 e339 ( .InEdge(Out21), .OutEdge(In80[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID340 e340 ( .InEdge(Out138), .OutEdge(In80[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID341 e341 ( .InEdge(Out413), .OutEdge(In80[6:6]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID81_INDEGREE1 n81 ( .InEdges(In81), .OutEdge(Out81),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID342 e342 ( .InEdge(Out258), .OutEdge(In81[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID82_INDEGREE1 n82 ( .InEdges(In82), .OutEdge(Out82),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID343 e343 ( .InEdge(Out448), .OutEdge(In82[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID83_INDEGREE6 n83 ( .InEdges(In83), .OutEdge(Out83),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID344 e344 ( .InEdge(Out479), .OutEdge(In83[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID345 e345 ( .InEdge(Out172), .OutEdge(In83[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID346 e346 ( .InEdge(Out8), .OutEdge(In83[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID347 e347 ( .InEdge(Out128), .OutEdge(In83[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID348 e348 ( .InEdge(Out108), .OutEdge(In83[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID349 e349 ( .InEdge(Out79), .OutEdge(In83[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID84_INDEGREE5 n84 ( .InEdges(In84), .OutEdge(Out84),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID350 e350 ( .InEdge(Out459), .OutEdge(In84[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID351 e351 ( .InEdge(Out443), .OutEdge(In84[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID352 e352 ( .InEdge(Out429), .OutEdge(In84[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID353 e353 ( .InEdge(Out290), .OutEdge(In84[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID354 e354 ( .InEdge(Out43), .OutEdge(In84[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID85_INDEGREE2 n85 ( .InEdges(In85), .OutEdge(Out85),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID355 e355 ( .InEdge(Out364), .OutEdge(In85[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID356 e356 ( .InEdge(Out507), .OutEdge(In85[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID86_INDEGREE1 n86 ( .InEdges(In86), .OutEdge(Out86),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID357 e357 ( .InEdge(Out204), .OutEdge(In86[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID87_INDEGREE3 n87 ( .InEdges(In87), .OutEdge(Out87),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID358 e358 ( .InEdge(Out207), .OutEdge(In87[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID359 e359 ( .InEdge(Out133), .OutEdge(In87[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID360 e360 ( .InEdge(Out231), .OutEdge(In87[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID88_INDEGREE5 n88 ( .InEdges(In88), .OutEdge(Out88),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID361 e361 ( .InEdge(Out180), .OutEdge(In88[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID362 e362 ( .InEdge(Out24), .OutEdge(In88[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID363 e363 ( .InEdge(Out265), .OutEdge(In88[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID364 e364 ( .InEdge(Out489), .OutEdge(In88[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID365 e365 ( .InEdge(Out423), .OutEdge(In88[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID89_INDEGREE7 n89 ( .InEdges(In89), .OutEdge(Out89),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID366 e366 ( .InEdge(Out235), .OutEdge(In89[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID367 e367 ( .InEdge(Out414), .OutEdge(In89[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID368 e368 ( .InEdge(Out6), .OutEdge(In89[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID369 e369 ( .InEdge(Out87), .OutEdge(In89[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID370 e370 ( .InEdge(Out149), .OutEdge(In89[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID371 e371 ( .InEdge(Out103), .OutEdge(In89[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID372 e372 ( .InEdge(Out399), .OutEdge(In89[6:6]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID90_INDEGREE3 n90 ( .InEdges(In90), .OutEdge(Out90),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID373 e373 ( .InEdge(Out340), .OutEdge(In90[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID374 e374 ( .InEdge(Out367), .OutEdge(In90[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID375 e375 ( .InEdge(Out392), .OutEdge(In90[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID91_INDEGREE6 n91 ( .InEdges(In91), .OutEdge(Out91),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID376 e376 ( .InEdge(Out246), .OutEdge(In91[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID377 e377 ( .InEdge(Out272), .OutEdge(In91[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID378 e378 ( .InEdge(Out302), .OutEdge(In91[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID379 e379 ( .InEdge(Out25), .OutEdge(In91[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID380 e380 ( .InEdge(Out380), .OutEdge(In91[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID381 e381 ( .InEdge(Out477), .OutEdge(In91[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID92_INDEGREE6 n92 ( .InEdges(In92), .OutEdge(Out92),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID382 e382 ( .InEdge(Out468), .OutEdge(In92[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID383 e383 ( .InEdge(Out483), .OutEdge(In92[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID384 e384 ( .InEdge(Out88), .OutEdge(In92[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID385 e385 ( .InEdge(Out497), .OutEdge(In92[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID386 e386 ( .InEdge(Out392), .OutEdge(In92[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID387 e387 ( .InEdge(Out350), .OutEdge(In92[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID93_INDEGREE3 n93 ( .InEdges(In93), .OutEdge(Out93),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID388 e388 ( .InEdge(Out452), .OutEdge(In93[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID389 e389 ( .InEdge(Out293), .OutEdge(In93[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID390 e390 ( .InEdge(Out61), .OutEdge(In93[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID94_INDEGREE1 n94 ( .InEdges(In94), .OutEdge(Out94),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID391 e391 ( .InEdge(Out350), .OutEdge(In94[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID95_INDEGREE6 n95 ( .InEdges(In95), .OutEdge(Out95),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID392 e392 ( .InEdge(Out431), .OutEdge(In95[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID393 e393 ( .InEdge(Out340), .OutEdge(In95[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID394 e394 ( .InEdge(Out246), .OutEdge(In95[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID395 e395 ( .InEdge(Out149), .OutEdge(In95[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID396 e396 ( .InEdge(Out18), .OutEdge(In95[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID397 e397 ( .InEdge(Out269), .OutEdge(In95[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID96_INDEGREE5 n96 ( .InEdges(In96), .OutEdge(Out96),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID398 e398 ( .InEdge(Out73), .OutEdge(In96[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID399 e399 ( .InEdge(Out16), .OutEdge(In96[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID400 e400 ( .InEdge(Out269), .OutEdge(In96[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID401 e401 ( .InEdge(Out364), .OutEdge(In96[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID402 e402 ( .InEdge(Out66), .OutEdge(In96[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID97_INDEGREE4 n97 ( .InEdges(In97), .OutEdge(Out97),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID403 e403 ( .InEdge(Out12), .OutEdge(In97[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID404 e404 ( .InEdge(Out21), .OutEdge(In97[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID405 e405 ( .InEdge(Out503), .OutEdge(In97[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID406 e406 ( .InEdge(Out49), .OutEdge(In97[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID98_INDEGREE6 n98 ( .InEdges(In98), .OutEdge(Out98),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID407 e407 ( .InEdge(Out97), .OutEdge(In98[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID408 e408 ( .InEdge(Out372), .OutEdge(In98[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID409 e409 ( .InEdge(Out401), .OutEdge(In98[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID410 e410 ( .InEdge(Out196), .OutEdge(In98[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID411 e411 ( .InEdge(Out420), .OutEdge(In98[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID412 e412 ( .InEdge(Out452), .OutEdge(In98[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID99_INDEGREE5 n99 ( .InEdges(In99), .OutEdge(Out99),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID413 e413 ( .InEdge(Out228), .OutEdge(In99[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID414 e414 ( .InEdge(Out488), .OutEdge(In99[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID415 e415 ( .InEdge(Out60), .OutEdge(In99[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID416 e416 ( .InEdge(Out185), .OutEdge(In99[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID417 e417 ( .InEdge(Out384), .OutEdge(In99[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID100_INDEGREE4 n100 ( .InEdges(In100), .OutEdge(Out100),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID418 e418 ( .InEdge(Out481), .OutEdge(In100[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID419 e419 ( .InEdge(Out202), .OutEdge(In100[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID420 e420 ( .InEdge(Out493), .OutEdge(In100[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID421 e421 ( .InEdge(Out113), .OutEdge(In100[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID101_INDEGREE4 n101 ( .InEdges(In101), .OutEdge(Out101),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID422 e422 ( .InEdge(Out311), .OutEdge(In101[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID423 e423 ( .InEdge(Out334), .OutEdge(In101[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID424 e424 ( .InEdge(Out57), .OutEdge(In101[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID425 e425 ( .InEdge(Out22), .OutEdge(In101[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID102_INDEGREE4 n102 ( .InEdges(In102), .OutEdge(Out102),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID426 e426 ( .InEdge(Out15), .OutEdge(In102[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID427 e427 ( .InEdge(Out409), .OutEdge(In102[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID428 e428 ( .InEdge(Out471), .OutEdge(In102[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID429 e429 ( .InEdge(Out48), .OutEdge(In102[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID103_INDEGREE3 n103 ( .InEdges(In103), .OutEdge(Out103),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID430 e430 ( .InEdge(Out23), .OutEdge(In103[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID431 e431 ( .InEdge(Out411), .OutEdge(In103[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID432 e432 ( .InEdge(Out360), .OutEdge(In103[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID104_INDEGREE5 n104 ( .InEdges(In104), .OutEdge(Out104),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID433 e433 ( .InEdge(Out121), .OutEdge(In104[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID434 e434 ( .InEdge(Out119), .OutEdge(In104[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID435 e435 ( .InEdge(Out128), .OutEdge(In104[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID436 e436 ( .InEdge(Out347), .OutEdge(In104[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID437 e437 ( .InEdge(Out367), .OutEdge(In104[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID105_INDEGREE3 n105 ( .InEdges(In105), .OutEdge(Out105),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID438 e438 ( .InEdge(Out493), .OutEdge(In105[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID439 e439 ( .InEdge(Out50), .OutEdge(In105[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID440 e440 ( .InEdge(Out380), .OutEdge(In105[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID106_INDEGREE7 n106 ( .InEdges(In106), .OutEdge(Out106),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID441 e441 ( .InEdge(Out116), .OutEdge(In106[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID442 e442 ( .InEdge(Out497), .OutEdge(In106[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID443 e443 ( .InEdge(Out304), .OutEdge(In106[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID444 e444 ( .InEdge(Out307), .OutEdge(In106[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID445 e445 ( .InEdge(Out415), .OutEdge(In106[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID446 e446 ( .InEdge(Out353), .OutEdge(In106[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID447 e447 ( .InEdge(Out41), .OutEdge(In106[6:6]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID107_INDEGREE5 n107 ( .InEdges(In107), .OutEdge(Out107),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID448 e448 ( .InEdge(Out211), .OutEdge(In107[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID449 e449 ( .InEdge(Out208), .OutEdge(In107[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID450 e450 ( .InEdge(Out263), .OutEdge(In107[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID451 e451 ( .InEdge(Out303), .OutEdge(In107[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID452 e452 ( .InEdge(Out5), .OutEdge(In107[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID108_INDEGREE5 n108 ( .InEdges(In108), .OutEdge(Out108),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID453 e453 ( .InEdge(Out63), .OutEdge(In108[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID454 e454 ( .InEdge(Out401), .OutEdge(In108[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID455 e455 ( .InEdge(Out104), .OutEdge(In108[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID456 e456 ( .InEdge(Out308), .OutEdge(In108[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID457 e457 ( .InEdge(Out499), .OutEdge(In108[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID109_INDEGREE2 n109 ( .InEdges(In109), .OutEdge(Out109),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID458 e458 ( .InEdge(Out225), .OutEdge(In109[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID459 e459 ( .InEdge(Out334), .OutEdge(In109[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID110_INDEGREE5 n110 ( .InEdges(In110), .OutEdge(Out110),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID460 e460 ( .InEdge(Out226), .OutEdge(In110[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID461 e461 ( .InEdge(Out17), .OutEdge(In110[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID462 e462 ( .InEdge(Out65), .OutEdge(In110[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID463 e463 ( .InEdge(Out56), .OutEdge(In110[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID464 e464 ( .InEdge(Out500), .OutEdge(In110[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID111_INDEGREE7 n111 ( .InEdges(In111), .OutEdge(Out111),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID465 e465 ( .InEdge(Out241), .OutEdge(In111[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID466 e466 ( .InEdge(Out281), .OutEdge(In111[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID467 e467 ( .InEdge(Out299), .OutEdge(In111[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID468 e468 ( .InEdge(Out428), .OutEdge(In111[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID469 e469 ( .InEdge(Out445), .OutEdge(In111[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID470 e470 ( .InEdge(Out398), .OutEdge(In111[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID471 e471 ( .InEdge(Out262), .OutEdge(In111[6:6]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID112_INDEGREE5 n112 ( .InEdges(In112), .OutEdge(Out112),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID472 e472 ( .InEdge(Out278), .OutEdge(In112[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID473 e473 ( .InEdge(Out69), .OutEdge(In112[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID474 e474 ( .InEdge(Out123), .OutEdge(In112[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID475 e475 ( .InEdge(Out25), .OutEdge(In112[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID476 e476 ( .InEdge(Out299), .OutEdge(In112[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID113_INDEGREE2 n113 ( .InEdges(In113), .OutEdge(Out113),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID477 e477 ( .InEdge(Out420), .OutEdge(In113[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID478 e478 ( .InEdge(Out413), .OutEdge(In113[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID114_INDEGREE3 n114 ( .InEdges(In114), .OutEdge(Out114),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID479 e479 ( .InEdge(Out52), .OutEdge(In114[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID480 e480 ( .InEdge(Out446), .OutEdge(In114[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID481 e481 ( .InEdge(Out424), .OutEdge(In114[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID115_INDEGREE4 n115 ( .InEdges(In115), .OutEdge(Out115),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID482 e482 ( .InEdge(Out196), .OutEdge(In115[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID483 e483 ( .InEdge(Out378), .OutEdge(In115[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID484 e484 ( .InEdge(Out468), .OutEdge(In115[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID485 e485 ( .InEdge(Out405), .OutEdge(In115[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID116_INDEGREE7 n116 ( .InEdges(In116), .OutEdge(Out116),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID486 e486 ( .InEdge(Out467), .OutEdge(In116[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID487 e487 ( .InEdge(Out362), .OutEdge(In116[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID488 e488 ( .InEdge(Out264), .OutEdge(In116[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID489 e489 ( .InEdge(Out169), .OutEdge(In116[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID490 e490 ( .InEdge(Out59), .OutEdge(In116[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID491 e491 ( .InEdge(Out420), .OutEdge(In116[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID492 e492 ( .InEdge(Out393), .OutEdge(In116[6:6]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID117_INDEGREE2 n117 ( .InEdges(In117), .OutEdge(Out117),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID493 e493 ( .InEdge(Out129), .OutEdge(In117[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID494 e494 ( .InEdge(Out172), .OutEdge(In117[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID118_INDEGREE2 n118 ( .InEdges(In118), .OutEdge(Out118),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID495 e495 ( .InEdge(Out486), .OutEdge(In118[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID496 e496 ( .InEdge(Out38), .OutEdge(In118[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID119_INDEGREE7 n119 ( .InEdges(In119), .OutEdge(Out119),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID497 e497 ( .InEdge(Out470), .OutEdge(In119[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID498 e498 ( .InEdge(Out202), .OutEdge(In119[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID499 e499 ( .InEdge(Out35), .OutEdge(In119[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID500 e500 ( .InEdge(Out203), .OutEdge(In119[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID501 e501 ( .InEdge(Out386), .OutEdge(In119[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID502 e502 ( .InEdge(Out306), .OutEdge(In119[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID503 e503 ( .InEdge(Out347), .OutEdge(In119[6:6]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID120_INDEGREE6 n120 ( .InEdges(In120), .OutEdge(Out120),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID504 e504 ( .InEdge(Out168), .OutEdge(In120[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID505 e505 ( .InEdge(Out68), .OutEdge(In120[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID506 e506 ( .InEdge(Out104), .OutEdge(In120[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID507 e507 ( .InEdge(Out263), .OutEdge(In120[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID508 e508 ( .InEdge(Out261), .OutEdge(In120[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID509 e509 ( .InEdge(Out45), .OutEdge(In120[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID121_INDEGREE6 n121 ( .InEdges(In121), .OutEdge(Out121),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID510 e510 ( .InEdge(Out303), .OutEdge(In121[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID511 e511 ( .InEdge(Out226), .OutEdge(In121[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID512 e512 ( .InEdge(Out407), .OutEdge(In121[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID513 e513 ( .InEdge(Out292), .OutEdge(In121[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID514 e514 ( .InEdge(Out225), .OutEdge(In121[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID515 e515 ( .InEdge(Out368), .OutEdge(In121[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID122_INDEGREE7 n122 ( .InEdges(In122), .OutEdge(Out122),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID516 e516 ( .InEdge(Out275), .OutEdge(In122[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID517 e517 ( .InEdge(Out62), .OutEdge(In122[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID518 e518 ( .InEdge(Out321), .OutEdge(In122[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID519 e519 ( .InEdge(Out408), .OutEdge(In122[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID520 e520 ( .InEdge(Out466), .OutEdge(In122[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID521 e521 ( .InEdge(Out45), .OutEdge(In122[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID522 e522 ( .InEdge(Out256), .OutEdge(In122[6:6]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID123_INDEGREE1 n123 ( .InEdges(In123), .OutEdge(Out123),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID523 e523 ( .InEdge(Out3), .OutEdge(In123[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID124_INDEGREE3 n124 ( .InEdges(In124), .OutEdge(Out124),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID524 e524 ( .InEdge(Out337), .OutEdge(In124[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID525 e525 ( .InEdge(Out284), .OutEdge(In124[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID526 e526 ( .InEdge(Out474), .OutEdge(In124[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID125_INDEGREE1 n125 ( .InEdges(In125), .OutEdge(Out125),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID527 e527 ( .InEdge(Out365), .OutEdge(In125[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID126_INDEGREE5 n126 ( .InEdges(In126), .OutEdge(Out126),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID528 e528 ( .InEdge(Out222), .OutEdge(In126[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID529 e529 ( .InEdge(Out431), .OutEdge(In126[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID530 e530 ( .InEdge(Out456), .OutEdge(In126[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID531 e531 ( .InEdge(Out507), .OutEdge(In126[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID532 e532 ( .InEdge(Out173), .OutEdge(In126[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID127_INDEGREE6 n127 ( .InEdges(In127), .OutEdge(Out127),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID533 e533 ( .InEdge(Out88), .OutEdge(In127[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID534 e534 ( .InEdge(Out456), .OutEdge(In127[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID535 e535 ( .InEdge(Out115), .OutEdge(In127[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID536 e536 ( .InEdge(Out271), .OutEdge(In127[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID537 e537 ( .InEdge(Out252), .OutEdge(In127[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID538 e538 ( .InEdge(Out385), .OutEdge(In127[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID128_INDEGREE3 n128 ( .InEdges(In128), .OutEdge(Out128),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID539 e539 ( .InEdge(Out173), .OutEdge(In128[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID540 e540 ( .InEdge(Out480), .OutEdge(In128[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID541 e541 ( .InEdge(Out239), .OutEdge(In128[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID129_INDEGREE3 n129 ( .InEdges(In129), .OutEdge(Out129),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID542 e542 ( .InEdge(Out128), .OutEdge(In129[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID543 e543 ( .InEdge(Out138), .OutEdge(In129[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID544 e544 ( .InEdge(Out242), .OutEdge(In129[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID130_INDEGREE2 n130 ( .InEdges(In130), .OutEdge(Out130),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID545 e545 ( .InEdge(Out359), .OutEdge(In130[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID546 e546 ( .InEdge(Out53), .OutEdge(In130[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID131_INDEGREE4 n131 ( .InEdges(In131), .OutEdge(Out131),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID547 e547 ( .InEdge(Out335), .OutEdge(In131[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID548 e548 ( .InEdge(Out435), .OutEdge(In131[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID549 e549 ( .InEdge(Out96), .OutEdge(In131[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID550 e550 ( .InEdge(Out367), .OutEdge(In131[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID132_INDEGREE5 n132 ( .InEdges(In132), .OutEdge(Out132),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID551 e551 ( .InEdge(Out342), .OutEdge(In132[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID552 e552 ( .InEdge(Out283), .OutEdge(In132[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID553 e553 ( .InEdge(Out203), .OutEdge(In132[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID554 e554 ( .InEdge(Out20), .OutEdge(In132[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID555 e555 ( .InEdge(Out116), .OutEdge(In132[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID133_INDEGREE7 n133 ( .InEdges(In133), .OutEdge(Out133),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID556 e556 ( .InEdge(Out94), .OutEdge(In133[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID557 e557 ( .InEdge(Out417), .OutEdge(In133[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID558 e558 ( .InEdge(Out451), .OutEdge(In133[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID559 e559 ( .InEdge(Out61), .OutEdge(In133[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID560 e560 ( .InEdge(Out291), .OutEdge(In133[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID561 e561 ( .InEdge(Out337), .OutEdge(In133[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID562 e562 ( .InEdge(Out195), .OutEdge(In133[6:6]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID134_INDEGREE3 n134 ( .InEdges(In134), .OutEdge(Out134),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID563 e563 ( .InEdge(Out17), .OutEdge(In134[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID564 e564 ( .InEdge(Out433), .OutEdge(In134[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID565 e565 ( .InEdge(Out280), .OutEdge(In134[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID135_INDEGREE7 n135 ( .InEdges(In135), .OutEdge(Out135),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID566 e566 ( .InEdge(Out73), .OutEdge(In135[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID567 e567 ( .InEdge(Out138), .OutEdge(In135[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID568 e568 ( .InEdge(Out213), .OutEdge(In135[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID569 e569 ( .InEdge(Out82), .OutEdge(In135[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID570 e570 ( .InEdge(Out289), .OutEdge(In135[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID571 e571 ( .InEdge(Out278), .OutEdge(In135[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID572 e572 ( .InEdge(Out444), .OutEdge(In135[6:6]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID136_INDEGREE5 n136 ( .InEdges(In136), .OutEdge(Out136),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID573 e573 ( .InEdge(Out403), .OutEdge(In136[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID574 e574 ( .InEdge(Out91), .OutEdge(In136[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID575 e575 ( .InEdge(Out110), .OutEdge(In136[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID576 e576 ( .InEdge(Out49), .OutEdge(In136[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID577 e577 ( .InEdge(Out229), .OutEdge(In136[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID137_INDEGREE3 n137 ( .InEdges(In137), .OutEdge(Out137),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID578 e578 ( .InEdge(Out485), .OutEdge(In137[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID579 e579 ( .InEdge(Out246), .OutEdge(In137[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID580 e580 ( .InEdge(Out158), .OutEdge(In137[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID138_INDEGREE1 n138 ( .InEdges(In138), .OutEdge(Out138),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID581 e581 ( .InEdge(Out279), .OutEdge(In138[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID139_INDEGREE2 n139 ( .InEdges(In139), .OutEdge(Out139),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID582 e582 ( .InEdge(Out436), .OutEdge(In139[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID583 e583 ( .InEdge(Out168), .OutEdge(In139[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID140_INDEGREE4 n140 ( .InEdges(In140), .OutEdge(Out140),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID584 e584 ( .InEdge(Out295), .OutEdge(In140[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID585 e585 ( .InEdge(Out127), .OutEdge(In140[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID586 e586 ( .InEdge(Out351), .OutEdge(In140[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID587 e587 ( .InEdge(Out306), .OutEdge(In140[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID141_INDEGREE7 n141 ( .InEdges(In141), .OutEdge(Out141),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID588 e588 ( .InEdge(Out95), .OutEdge(In141[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID589 e589 ( .InEdge(Out242), .OutEdge(In141[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID590 e590 ( .InEdge(Out379), .OutEdge(In141[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID591 e591 ( .InEdge(Out175), .OutEdge(In141[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID592 e592 ( .InEdge(Out263), .OutEdge(In141[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID593 e593 ( .InEdge(Out487), .OutEdge(In141[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID594 e594 ( .InEdge(Out140), .OutEdge(In141[6:6]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID142_INDEGREE1 n142 ( .InEdges(In142), .OutEdge(Out142),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID595 e595 ( .InEdge(Out255), .OutEdge(In142[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID143_INDEGREE6 n143 ( .InEdges(In143), .OutEdge(Out143),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID596 e596 ( .InEdge(Out160), .OutEdge(In143[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID597 e597 ( .InEdge(Out496), .OutEdge(In143[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID598 e598 ( .InEdge(Out430), .OutEdge(In143[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID599 e599 ( .InEdge(Out354), .OutEdge(In143[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID600 e600 ( .InEdge(Out309), .OutEdge(In143[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID601 e601 ( .InEdge(Out133), .OutEdge(In143[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID144_INDEGREE6 n144 ( .InEdges(In144), .OutEdge(Out144),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID602 e602 ( .InEdge(Out15), .OutEdge(In144[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID603 e603 ( .InEdge(Out265), .OutEdge(In144[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID604 e604 ( .InEdge(Out256), .OutEdge(In144[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID605 e605 ( .InEdge(Out169), .OutEdge(In144[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID606 e606 ( .InEdge(Out402), .OutEdge(In144[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID607 e607 ( .InEdge(Out314), .OutEdge(In144[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID145_INDEGREE3 n145 ( .InEdges(In145), .OutEdge(Out145),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID608 e608 ( .InEdge(Out499), .OutEdge(In145[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID609 e609 ( .InEdge(Out0), .OutEdge(In145[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID610 e610 ( .InEdge(Out286), .OutEdge(In145[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID146_INDEGREE3 n146 ( .InEdges(In146), .OutEdge(Out146),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID611 e611 ( .InEdge(Out30), .OutEdge(In146[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID612 e612 ( .InEdge(Out230), .OutEdge(In146[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID613 e613 ( .InEdge(Out106), .OutEdge(In146[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID147_INDEGREE5 n147 ( .InEdges(In147), .OutEdge(Out147),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID614 e614 ( .InEdge(Out308), .OutEdge(In147[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID615 e615 ( .InEdge(Out7), .OutEdge(In147[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID616 e616 ( .InEdge(Out359), .OutEdge(In147[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID617 e617 ( .InEdge(Out333), .OutEdge(In147[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID618 e618 ( .InEdge(Out477), .OutEdge(In147[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID148_INDEGREE7 n148 ( .InEdges(In148), .OutEdge(Out148),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID619 e619 ( .InEdge(Out340), .OutEdge(In148[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID620 e620 ( .InEdge(Out395), .OutEdge(In148[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID621 e621 ( .InEdge(Out184), .OutEdge(In148[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID622 e622 ( .InEdge(Out256), .OutEdge(In148[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID623 e623 ( .InEdge(Out161), .OutEdge(In148[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID624 e624 ( .InEdge(Out183), .OutEdge(In148[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID625 e625 ( .InEdge(Out309), .OutEdge(In148[6:6]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID149_INDEGREE4 n149 ( .InEdges(In149), .OutEdge(Out149),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID626 e626 ( .InEdge(Out157), .OutEdge(In149[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID627 e627 ( .InEdge(Out500), .OutEdge(In149[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID628 e628 ( .InEdge(Out165), .OutEdge(In149[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID629 e629 ( .InEdge(Out187), .OutEdge(In149[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID150_INDEGREE6 n150 ( .InEdges(In150), .OutEdge(Out150),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID630 e630 ( .InEdge(Out1), .OutEdge(In150[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID631 e631 ( .InEdge(Out54), .OutEdge(In150[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID632 e632 ( .InEdge(Out172), .OutEdge(In150[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID633 e633 ( .InEdge(Out409), .OutEdge(In150[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID634 e634 ( .InEdge(Out378), .OutEdge(In150[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID635 e635 ( .InEdge(Out268), .OutEdge(In150[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID151_INDEGREE3 n151 ( .InEdges(In151), .OutEdge(Out151),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID636 e636 ( .InEdge(Out254), .OutEdge(In151[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID637 e637 ( .InEdge(Out257), .OutEdge(In151[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID638 e638 ( .InEdge(Out367), .OutEdge(In151[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID152_INDEGREE7 n152 ( .InEdges(In152), .OutEdge(Out152),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID639 e639 ( .InEdge(Out266), .OutEdge(In152[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID640 e640 ( .InEdge(Out499), .OutEdge(In152[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID641 e641 ( .InEdge(Out157), .OutEdge(In152[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID642 e642 ( .InEdge(Out350), .OutEdge(In152[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID643 e643 ( .InEdge(Out129), .OutEdge(In152[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID644 e644 ( .InEdge(Out352), .OutEdge(In152[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID645 e645 ( .InEdge(Out102), .OutEdge(In152[6:6]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID153_INDEGREE4 n153 ( .InEdges(In153), .OutEdge(Out153),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID646 e646 ( .InEdge(Out116), .OutEdge(In153[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID647 e647 ( .InEdge(Out237), .OutEdge(In153[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID648 e648 ( .InEdge(Out287), .OutEdge(In153[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID649 e649 ( .InEdge(Out283), .OutEdge(In153[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID154_INDEGREE7 n154 ( .InEdges(In154), .OutEdge(Out154),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID650 e650 ( .InEdge(Out446), .OutEdge(In154[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID651 e651 ( .InEdge(Out256), .OutEdge(In154[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID652 e652 ( .InEdge(Out193), .OutEdge(In154[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID653 e653 ( .InEdge(Out149), .OutEdge(In154[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID654 e654 ( .InEdge(Out424), .OutEdge(In154[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID655 e655 ( .InEdge(Out278), .OutEdge(In154[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID656 e656 ( .InEdge(Out249), .OutEdge(In154[6:6]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID155_INDEGREE1 n155 ( .InEdges(In155), .OutEdge(Out155),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID657 e657 ( .InEdge(Out372), .OutEdge(In155[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID156_INDEGREE5 n156 ( .InEdges(In156), .OutEdge(Out156),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID658 e658 ( .InEdge(Out94), .OutEdge(In156[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID659 e659 ( .InEdge(Out392), .OutEdge(In156[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID660 e660 ( .InEdge(Out315), .OutEdge(In156[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID661 e661 ( .InEdge(Out394), .OutEdge(In156[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID662 e662 ( .InEdge(Out354), .OutEdge(In156[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID157_INDEGREE7 n157 ( .InEdges(In157), .OutEdge(Out157),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID663 e663 ( .InEdge(Out168), .OutEdge(In157[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID664 e664 ( .InEdge(Out412), .OutEdge(In157[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID665 e665 ( .InEdge(Out18), .OutEdge(In157[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID666 e666 ( .InEdge(Out45), .OutEdge(In157[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID667 e667 ( .InEdge(Out162), .OutEdge(In157[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID668 e668 ( .InEdge(Out464), .OutEdge(In157[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID669 e669 ( .InEdge(Out4), .OutEdge(In157[6:6]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID158_INDEGREE2 n158 ( .InEdges(In158), .OutEdge(Out158),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID670 e670 ( .InEdge(Out384), .OutEdge(In158[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID671 e671 ( .InEdge(Out117), .OutEdge(In158[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID159_INDEGREE7 n159 ( .InEdges(In159), .OutEdge(Out159),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID672 e672 ( .InEdge(Out262), .OutEdge(In159[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID673 e673 ( .InEdge(Out49), .OutEdge(In159[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID674 e674 ( .InEdge(Out18), .OutEdge(In159[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID675 e675 ( .InEdge(Out288), .OutEdge(In159[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID676 e676 ( .InEdge(Out363), .OutEdge(In159[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID677 e677 ( .InEdge(Out90), .OutEdge(In159[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID678 e678 ( .InEdge(Out74), .OutEdge(In159[6:6]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID160_INDEGREE7 n160 ( .InEdges(In160), .OutEdge(Out160),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID679 e679 ( .InEdge(Out99), .OutEdge(In160[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID680 e680 ( .InEdge(Out297), .OutEdge(In160[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID681 e681 ( .InEdge(Out118), .OutEdge(In160[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID682 e682 ( .InEdge(Out48), .OutEdge(In160[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID683 e683 ( .InEdge(Out166), .OutEdge(In160[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID684 e684 ( .InEdge(Out403), .OutEdge(In160[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID685 e685 ( .InEdge(Out372), .OutEdge(In160[6:6]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID161_INDEGREE4 n161 ( .InEdges(In161), .OutEdge(Out161),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID686 e686 ( .InEdge(Out334), .OutEdge(In161[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID687 e687 ( .InEdge(Out53), .OutEdge(In161[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID688 e688 ( .InEdge(Out287), .OutEdge(In161[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID689 e689 ( .InEdge(Out81), .OutEdge(In161[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID162_INDEGREE2 n162 ( .InEdges(In162), .OutEdge(Out162),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID690 e690 ( .InEdge(Out500), .OutEdge(In162[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID691 e691 ( .InEdge(Out385), .OutEdge(In162[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID163_INDEGREE7 n163 ( .InEdges(In163), .OutEdge(Out163),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID692 e692 ( .InEdge(Out408), .OutEdge(In163[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID693 e693 ( .InEdge(Out41), .OutEdge(In163[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID694 e694 ( .InEdge(Out189), .OutEdge(In163[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID695 e695 ( .InEdge(Out268), .OutEdge(In163[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID696 e696 ( .InEdge(Out479), .OutEdge(In163[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID697 e697 ( .InEdge(Out261), .OutEdge(In163[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID698 e698 ( .InEdge(Out504), .OutEdge(In163[6:6]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID164_INDEGREE5 n164 ( .InEdges(In164), .OutEdge(Out164),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID699 e699 ( .InEdge(Out509), .OutEdge(In164[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID700 e700 ( .InEdge(Out302), .OutEdge(In164[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID701 e701 ( .InEdge(Out149), .OutEdge(In164[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID702 e702 ( .InEdge(Out77), .OutEdge(In164[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID703 e703 ( .InEdge(Out487), .OutEdge(In164[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID165_INDEGREE1 n165 ( .InEdges(In165), .OutEdge(Out165),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID704 e704 ( .InEdge(Out357), .OutEdge(In165[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID166_INDEGREE1 n166 ( .InEdges(In166), .OutEdge(Out166),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID705 e705 ( .InEdge(Out182), .OutEdge(In166[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID167_INDEGREE6 n167 ( .InEdges(In167), .OutEdge(Out167),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID706 e706 ( .InEdge(Out36), .OutEdge(In167[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID707 e707 ( .InEdge(Out384), .OutEdge(In167[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID708 e708 ( .InEdge(Out391), .OutEdge(In167[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID709 e709 ( .InEdge(Out323), .OutEdge(In167[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID710 e710 ( .InEdge(Out18), .OutEdge(In167[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID711 e711 ( .InEdge(Out237), .OutEdge(In167[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID168_INDEGREE1 n168 ( .InEdges(In168), .OutEdge(Out168),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID712 e712 ( .InEdge(Out435), .OutEdge(In168[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID169_INDEGREE4 n169 ( .InEdges(In169), .OutEdge(Out169),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID713 e713 ( .InEdge(Out214), .OutEdge(In169[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID714 e714 ( .InEdge(Out246), .OutEdge(In169[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID715 e715 ( .InEdge(Out69), .OutEdge(In169[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID716 e716 ( .InEdge(Out49), .OutEdge(In169[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID170_INDEGREE5 n170 ( .InEdges(In170), .OutEdge(Out170),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID717 e717 ( .InEdge(Out189), .OutEdge(In170[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID718 e718 ( .InEdge(Out468), .OutEdge(In170[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID719 e719 ( .InEdge(Out238), .OutEdge(In170[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID720 e720 ( .InEdge(Out21), .OutEdge(In170[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID721 e721 ( .InEdge(Out445), .OutEdge(In170[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID171_INDEGREE5 n171 ( .InEdges(In171), .OutEdge(Out171),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID722 e722 ( .InEdge(Out268), .OutEdge(In171[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID723 e723 ( .InEdge(Out139), .OutEdge(In171[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID724 e724 ( .InEdge(Out287), .OutEdge(In171[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID725 e725 ( .InEdge(Out406), .OutEdge(In171[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID726 e726 ( .InEdge(Out35), .OutEdge(In171[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID172_INDEGREE7 n172 ( .InEdges(In172), .OutEdge(Out172),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID727 e727 ( .InEdge(Out237), .OutEdge(In172[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID728 e728 ( .InEdge(Out294), .OutEdge(In172[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID729 e729 ( .InEdge(Out216), .OutEdge(In172[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID730 e730 ( .InEdge(Out258), .OutEdge(In172[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID731 e731 ( .InEdge(Out316), .OutEdge(In172[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID732 e732 ( .InEdge(Out239), .OutEdge(In172[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID733 e733 ( .InEdge(Out245), .OutEdge(In172[6:6]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID173_INDEGREE2 n173 ( .InEdges(In173), .OutEdge(Out173),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID734 e734 ( .InEdge(Out208), .OutEdge(In173[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID735 e735 ( .InEdge(Out292), .OutEdge(In173[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID174_INDEGREE2 n174 ( .InEdges(In174), .OutEdge(Out174),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID736 e736 ( .InEdge(Out501), .OutEdge(In174[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID737 e737 ( .InEdge(Out308), .OutEdge(In174[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID175_INDEGREE1 n175 ( .InEdges(In175), .OutEdge(Out175),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID738 e738 ( .InEdge(Out224), .OutEdge(In175[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID176_INDEGREE5 n176 ( .InEdges(In176), .OutEdge(Out176),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID739 e739 ( .InEdge(Out268), .OutEdge(In176[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID740 e740 ( .InEdge(Out430), .OutEdge(In176[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID741 e741 ( .InEdge(Out8), .OutEdge(In176[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID742 e742 ( .InEdge(Out269), .OutEdge(In176[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID743 e743 ( .InEdge(Out243), .OutEdge(In176[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID177_INDEGREE1 n177 ( .InEdges(In177), .OutEdge(Out177),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID744 e744 ( .InEdge(Out265), .OutEdge(In177[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID178_INDEGREE5 n178 ( .InEdges(In178), .OutEdge(Out178),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID745 e745 ( .InEdge(Out163), .OutEdge(In178[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID746 e746 ( .InEdge(Out274), .OutEdge(In178[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID747 e747 ( .InEdge(Out126), .OutEdge(In178[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID748 e748 ( .InEdge(Out228), .OutEdge(In178[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID749 e749 ( .InEdge(Out22), .OutEdge(In178[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID179_INDEGREE7 n179 ( .InEdges(In179), .OutEdge(Out179),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID750 e750 ( .InEdge(Out194), .OutEdge(In179[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID751 e751 ( .InEdge(Out250), .OutEdge(In179[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID752 e752 ( .InEdge(Out140), .OutEdge(In179[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID753 e753 ( .InEdge(Out40), .OutEdge(In179[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID754 e754 ( .InEdge(Out343), .OutEdge(In179[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID755 e755 ( .InEdge(Out81), .OutEdge(In179[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID756 e756 ( .InEdge(Out504), .OutEdge(In179[6:6]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID180_INDEGREE6 n180 ( .InEdges(In180), .OutEdge(Out180),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID757 e757 ( .InEdge(Out419), .OutEdge(In180[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID758 e758 ( .InEdge(Out190), .OutEdge(In180[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID759 e759 ( .InEdge(Out285), .OutEdge(In180[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID760 e760 ( .InEdge(Out297), .OutEdge(In180[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID761 e761 ( .InEdge(Out343), .OutEdge(In180[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID762 e762 ( .InEdge(Out222), .OutEdge(In180[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID181_INDEGREE7 n181 ( .InEdges(In181), .OutEdge(Out181),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID763 e763 ( .InEdge(Out219), .OutEdge(In181[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID764 e764 ( .InEdge(Out210), .OutEdge(In181[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID765 e765 ( .InEdge(Out124), .OutEdge(In181[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID766 e766 ( .InEdge(Out447), .OutEdge(In181[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID767 e767 ( .InEdge(Out173), .OutEdge(In181[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID768 e768 ( .InEdge(Out288), .OutEdge(In181[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID769 e769 ( .InEdge(Out106), .OutEdge(In181[6:6]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID182_INDEGREE7 n182 ( .InEdges(In182), .OutEdge(Out182),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID770 e770 ( .InEdge(Out434), .OutEdge(In182[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID771 e771 ( .InEdge(Out362), .OutEdge(In182[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID772 e772 ( .InEdge(Out201), .OutEdge(In182[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID773 e773 ( .InEdge(Out62), .OutEdge(In182[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID774 e774 ( .InEdge(Out461), .OutEdge(In182[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID775 e775 ( .InEdge(Out88), .OutEdge(In182[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID776 e776 ( .InEdge(Out21), .OutEdge(In182[6:6]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID183_INDEGREE4 n183 ( .InEdges(In183), .OutEdge(Out183),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID777 e777 ( .InEdge(Out379), .OutEdge(In183[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID778 e778 ( .InEdge(Out124), .OutEdge(In183[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID779 e779 ( .InEdge(Out294), .OutEdge(In183[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID780 e780 ( .InEdge(Out433), .OutEdge(In183[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID184_INDEGREE7 n184 ( .InEdges(In184), .OutEdge(Out184),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID781 e781 ( .InEdge(Out205), .OutEdge(In184[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID782 e782 ( .InEdge(Out413), .OutEdge(In184[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID783 e783 ( .InEdge(Out5), .OutEdge(In184[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID784 e784 ( .InEdge(Out111), .OutEdge(In184[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID785 e785 ( .InEdge(Out355), .OutEdge(In184[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID786 e786 ( .InEdge(Out6), .OutEdge(In184[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID787 e787 ( .InEdge(Out318), .OutEdge(In184[6:6]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID185_INDEGREE1 n185 ( .InEdges(In185), .OutEdge(Out185),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID788 e788 ( .InEdge(Out359), .OutEdge(In185[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID186_INDEGREE1 n186 ( .InEdges(In186), .OutEdge(Out186),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID789 e789 ( .InEdge(Out326), .OutEdge(In186[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID187_INDEGREE3 n187 ( .InEdges(In187), .OutEdge(Out187),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID790 e790 ( .InEdge(Out57), .OutEdge(In187[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID791 e791 ( .InEdge(Out423), .OutEdge(In187[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID792 e792 ( .InEdge(Out237), .OutEdge(In187[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID188_INDEGREE5 n188 ( .InEdges(In188), .OutEdge(Out188),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID793 e793 ( .InEdge(Out337), .OutEdge(In188[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID794 e794 ( .InEdge(Out11), .OutEdge(In188[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID795 e795 ( .InEdge(Out328), .OutEdge(In188[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID796 e796 ( .InEdge(Out356), .OutEdge(In188[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID797 e797 ( .InEdge(Out380), .OutEdge(In188[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID189_INDEGREE7 n189 ( .InEdges(In189), .OutEdge(Out189),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID798 e798 ( .InEdge(Out84), .OutEdge(In189[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID799 e799 ( .InEdge(Out447), .OutEdge(In189[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID800 e800 ( .InEdge(Out449), .OutEdge(In189[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID801 e801 ( .InEdge(Out402), .OutEdge(In189[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID802 e802 ( .InEdge(Out301), .OutEdge(In189[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID803 e803 ( .InEdge(Out37), .OutEdge(In189[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID804 e804 ( .InEdge(Out389), .OutEdge(In189[6:6]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID190_INDEGREE7 n190 ( .InEdges(In190), .OutEdge(Out190),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID805 e805 ( .InEdge(Out279), .OutEdge(In190[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID806 e806 ( .InEdge(Out371), .OutEdge(In190[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID807 e807 ( .InEdge(Out372), .OutEdge(In190[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID808 e808 ( .InEdge(Out139), .OutEdge(In190[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID809 e809 ( .InEdge(Out232), .OutEdge(In190[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID810 e810 ( .InEdge(Out339), .OutEdge(In190[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID811 e811 ( .InEdge(Out120), .OutEdge(In190[6:6]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID191_INDEGREE2 n191 ( .InEdges(In191), .OutEdge(Out191),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID812 e812 ( .InEdge(Out144), .OutEdge(In191[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID813 e813 ( .InEdge(Out3), .OutEdge(In191[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID192_INDEGREE6 n192 ( .InEdges(In192), .OutEdge(Out192),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID814 e814 ( .InEdge(Out184), .OutEdge(In192[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID815 e815 ( .InEdge(Out240), .OutEdge(In192[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID816 e816 ( .InEdge(Out435), .OutEdge(In192[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID817 e817 ( .InEdge(Out233), .OutEdge(In192[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID818 e818 ( .InEdge(Out124), .OutEdge(In192[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID819 e819 ( .InEdge(Out417), .OutEdge(In192[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID193_INDEGREE6 n193 ( .InEdges(In193), .OutEdge(Out193),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID820 e820 ( .InEdge(Out66), .OutEdge(In193[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID821 e821 ( .InEdge(Out231), .OutEdge(In193[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID822 e822 ( .InEdge(Out82), .OutEdge(In193[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID823 e823 ( .InEdge(Out355), .OutEdge(In193[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID824 e824 ( .InEdge(Out236), .OutEdge(In193[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID825 e825 ( .InEdge(Out485), .OutEdge(In193[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID194_INDEGREE1 n194 ( .InEdges(In194), .OutEdge(Out194),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID826 e826 ( .InEdge(Out346), .OutEdge(In194[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID195_INDEGREE3 n195 ( .InEdges(In195), .OutEdge(Out195),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID827 e827 ( .InEdge(Out375), .OutEdge(In195[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID828 e828 ( .InEdge(Out21), .OutEdge(In195[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID829 e829 ( .InEdge(Out336), .OutEdge(In195[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID196_INDEGREE5 n196 ( .InEdges(In196), .OutEdge(Out196),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID830 e830 ( .InEdge(Out439), .OutEdge(In196[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID831 e831 ( .InEdge(Out346), .OutEdge(In196[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID832 e832 ( .InEdge(Out348), .OutEdge(In196[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID833 e833 ( .InEdge(Out226), .OutEdge(In196[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID834 e834 ( .InEdge(Out10), .OutEdge(In196[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID197_INDEGREE3 n197 ( .InEdges(In197), .OutEdge(Out197),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID835 e835 ( .InEdge(Out106), .OutEdge(In197[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID836 e836 ( .InEdge(Out79), .OutEdge(In197[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID837 e837 ( .InEdge(Out349), .OutEdge(In197[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID198_INDEGREE3 n198 ( .InEdges(In198), .OutEdge(Out198),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID838 e838 ( .InEdge(Out78), .OutEdge(In198[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID839 e839 ( .InEdge(Out377), .OutEdge(In198[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID840 e840 ( .InEdge(Out269), .OutEdge(In198[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID199_INDEGREE7 n199 ( .InEdges(In199), .OutEdge(Out199),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID841 e841 ( .InEdge(Out409), .OutEdge(In199[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID842 e842 ( .InEdge(Out503), .OutEdge(In199[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID843 e843 ( .InEdge(Out339), .OutEdge(In199[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID844 e844 ( .InEdge(Out260), .OutEdge(In199[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID845 e845 ( .InEdge(Out120), .OutEdge(In199[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID846 e846 ( .InEdge(Out476), .OutEdge(In199[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID847 e847 ( .InEdge(Out133), .OutEdge(In199[6:6]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID200_INDEGREE1 n200 ( .InEdges(In200), .OutEdge(Out200),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID848 e848 ( .InEdge(Out487), .OutEdge(In200[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID201_INDEGREE2 n201 ( .InEdges(In201), .OutEdge(Out201),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID849 e849 ( .InEdge(Out190), .OutEdge(In201[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID850 e850 ( .InEdge(Out309), .OutEdge(In201[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID202_INDEGREE5 n202 ( .InEdges(In202), .OutEdge(Out202),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID851 e851 ( .InEdge(Out461), .OutEdge(In202[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID852 e852 ( .InEdge(Out429), .OutEdge(In202[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID853 e853 ( .InEdge(Out72), .OutEdge(In202[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID854 e854 ( .InEdge(Out176), .OutEdge(In202[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID855 e855 ( .InEdge(Out329), .OutEdge(In202[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID203_INDEGREE3 n203 ( .InEdges(In203), .OutEdge(Out203),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID856 e856 ( .InEdge(Out323), .OutEdge(In203[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID857 e857 ( .InEdge(Out282), .OutEdge(In203[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID858 e858 ( .InEdge(Out320), .OutEdge(In203[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID204_INDEGREE6 n204 ( .InEdges(In204), .OutEdge(Out204),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID859 e859 ( .InEdge(Out276), .OutEdge(In204[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID860 e860 ( .InEdge(Out394), .OutEdge(In204[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID861 e861 ( .InEdge(Out329), .OutEdge(In204[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID862 e862 ( .InEdge(Out249), .OutEdge(In204[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID863 e863 ( .InEdge(Out494), .OutEdge(In204[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID864 e864 ( .InEdge(Out192), .OutEdge(In204[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID205_INDEGREE3 n205 ( .InEdges(In205), .OutEdge(Out205),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID865 e865 ( .InEdge(Out285), .OutEdge(In205[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID866 e866 ( .InEdge(Out222), .OutEdge(In205[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID867 e867 ( .InEdge(Out295), .OutEdge(In205[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID206_INDEGREE3 n206 ( .InEdges(In206), .OutEdge(Out206),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID868 e868 ( .InEdge(Out82), .OutEdge(In206[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID869 e869 ( .InEdge(Out391), .OutEdge(In206[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID870 e870 ( .InEdge(Out475), .OutEdge(In206[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID207_INDEGREE2 n207 ( .InEdges(In207), .OutEdge(Out207),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID871 e871 ( .InEdge(Out403), .OutEdge(In207[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID872 e872 ( .InEdge(Out12), .OutEdge(In207[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID208_INDEGREE5 n208 ( .InEdges(In208), .OutEdge(Out208),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID873 e873 ( .InEdge(Out148), .OutEdge(In208[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID874 e874 ( .InEdge(Out432), .OutEdge(In208[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID875 e875 ( .InEdge(Out301), .OutEdge(In208[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID876 e876 ( .InEdge(Out415), .OutEdge(In208[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID877 e877 ( .InEdge(Out134), .OutEdge(In208[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID209_INDEGREE2 n209 ( .InEdges(In209), .OutEdge(Out209),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID878 e878 ( .InEdge(Out463), .OutEdge(In209[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID879 e879 ( .InEdge(Out43), .OutEdge(In209[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID210_INDEGREE6 n210 ( .InEdges(In210), .OutEdge(Out210),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID880 e880 ( .InEdge(Out479), .OutEdge(In210[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID881 e881 ( .InEdge(Out450), .OutEdge(In210[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID882 e882 ( .InEdge(Out335), .OutEdge(In210[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID883 e883 ( .InEdge(Out249), .OutEdge(In210[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID884 e884 ( .InEdge(Out207), .OutEdge(In210[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID885 e885 ( .InEdge(Out306), .OutEdge(In210[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID211_INDEGREE6 n211 ( .InEdges(In211), .OutEdge(Out211),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID886 e886 ( .InEdge(Out378), .OutEdge(In211[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID887 e887 ( .InEdge(Out418), .OutEdge(In211[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID888 e888 ( .InEdge(Out55), .OutEdge(In211[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID889 e889 ( .InEdge(Out340), .OutEdge(In211[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID890 e890 ( .InEdge(Out375), .OutEdge(In211[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID891 e891 ( .InEdge(Out92), .OutEdge(In211[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID212_INDEGREE2 n212 ( .InEdges(In212), .OutEdge(Out212),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID892 e892 ( .InEdge(Out145), .OutEdge(In212[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID893 e893 ( .InEdge(Out413), .OutEdge(In212[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID213_INDEGREE2 n213 ( .InEdges(In213), .OutEdge(Out213),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID894 e894 ( .InEdge(Out227), .OutEdge(In213[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID895 e895 ( .InEdge(Out165), .OutEdge(In213[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID214_INDEGREE7 n214 ( .InEdges(In214), .OutEdge(Out214),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID896 e896 ( .InEdge(Out237), .OutEdge(In214[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID897 e897 ( .InEdge(Out143), .OutEdge(In214[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID898 e898 ( .InEdge(Out23), .OutEdge(In214[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID899 e899 ( .InEdge(Out69), .OutEdge(In214[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID900 e900 ( .InEdge(Out380), .OutEdge(In214[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID901 e901 ( .InEdge(Out222), .OutEdge(In214[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID902 e902 ( .InEdge(Out4), .OutEdge(In214[6:6]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID215_INDEGREE1 n215 ( .InEdges(In215), .OutEdge(Out215),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID903 e903 ( .InEdge(Out52), .OutEdge(In215[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID216_INDEGREE6 n216 ( .InEdges(In216), .OutEdge(Out216),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID904 e904 ( .InEdge(Out332), .OutEdge(In216[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID905 e905 ( .InEdge(Out115), .OutEdge(In216[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID906 e906 ( .InEdge(Out348), .OutEdge(In216[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID907 e907 ( .InEdge(Out176), .OutEdge(In216[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID908 e908 ( .InEdge(Out393), .OutEdge(In216[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID909 e909 ( .InEdge(Out369), .OutEdge(In216[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID217_INDEGREE4 n217 ( .InEdges(In217), .OutEdge(Out217),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID910 e910 ( .InEdge(Out457), .OutEdge(In217[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID911 e911 ( .InEdge(Out362), .OutEdge(In217[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID912 e912 ( .InEdge(Out165), .OutEdge(In217[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID913 e913 ( .InEdge(Out481), .OutEdge(In217[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID218_INDEGREE2 n218 ( .InEdges(In218), .OutEdge(Out218),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID914 e914 ( .InEdge(Out421), .OutEdge(In218[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID915 e915 ( .InEdge(Out62), .OutEdge(In218[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID219_INDEGREE3 n219 ( .InEdges(In219), .OutEdge(Out219),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID916 e916 ( .InEdge(Out115), .OutEdge(In219[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID917 e917 ( .InEdge(Out120), .OutEdge(In219[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID918 e918 ( .InEdge(Out334), .OutEdge(In219[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID220_INDEGREE5 n220 ( .InEdges(In220), .OutEdge(Out220),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID919 e919 ( .InEdge(Out11), .OutEdge(In220[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID920 e920 ( .InEdge(Out449), .OutEdge(In220[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID921 e921 ( .InEdge(Out158), .OutEdge(In220[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID922 e922 ( .InEdge(Out250), .OutEdge(In220[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID923 e923 ( .InEdge(Out151), .OutEdge(In220[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID221_INDEGREE3 n221 ( .InEdges(In221), .OutEdge(Out221),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID924 e924 ( .InEdge(Out209), .OutEdge(In221[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID925 e925 ( .InEdge(Out435), .OutEdge(In221[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID926 e926 ( .InEdge(Out323), .OutEdge(In221[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID222_INDEGREE1 n222 ( .InEdges(In222), .OutEdge(Out222),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID927 e927 ( .InEdge(Out479), .OutEdge(In222[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID223_INDEGREE3 n223 ( .InEdges(In223), .OutEdge(Out223),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID928 e928 ( .InEdge(Out365), .OutEdge(In223[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID929 e929 ( .InEdge(Out362), .OutEdge(In223[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID930 e930 ( .InEdge(Out389), .OutEdge(In223[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID224_INDEGREE7 n224 ( .InEdges(In224), .OutEdge(Out224),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID931 e931 ( .InEdge(Out499), .OutEdge(In224[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID932 e932 ( .InEdge(Out261), .OutEdge(In224[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID933 e933 ( .InEdge(Out490), .OutEdge(In224[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID934 e934 ( .InEdge(Out283), .OutEdge(In224[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID935 e935 ( .InEdge(Out432), .OutEdge(In224[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID936 e936 ( .InEdge(Out360), .OutEdge(In224[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID937 e937 ( .InEdge(Out154), .OutEdge(In224[6:6]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID225_INDEGREE5 n225 ( .InEdges(In225), .OutEdge(Out225),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID938 e938 ( .InEdge(Out237), .OutEdge(In225[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID939 e939 ( .InEdge(Out339), .OutEdge(In225[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID940 e940 ( .InEdge(Out335), .OutEdge(In225[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID941 e941 ( .InEdge(Out207), .OutEdge(In225[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID942 e942 ( .InEdge(Out62), .OutEdge(In225[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID226_INDEGREE5 n226 ( .InEdges(In226), .OutEdge(Out226),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID943 e943 ( .InEdge(Out443), .OutEdge(In226[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID944 e944 ( .InEdge(Out20), .OutEdge(In226[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID945 e945 ( .InEdge(Out27), .OutEdge(In226[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID946 e946 ( .InEdge(Out17), .OutEdge(In226[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID947 e947 ( .InEdge(Out314), .OutEdge(In226[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID227_INDEGREE1 n227 ( .InEdges(In227), .OutEdge(Out227),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID948 e948 ( .InEdge(Out11), .OutEdge(In227[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID228_INDEGREE2 n228 ( .InEdges(In228), .OutEdge(Out228),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID949 e949 ( .InEdge(Out29), .OutEdge(In228[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID950 e950 ( .InEdge(Out225), .OutEdge(In228[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID229_INDEGREE6 n229 ( .InEdges(In229), .OutEdge(Out229),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID951 e951 ( .InEdge(Out470), .OutEdge(In229[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID952 e952 ( .InEdge(Out344), .OutEdge(In229[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID953 e953 ( .InEdge(Out16), .OutEdge(In229[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID954 e954 ( .InEdge(Out215), .OutEdge(In229[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID955 e955 ( .InEdge(Out56), .OutEdge(In229[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID956 e956 ( .InEdge(Out61), .OutEdge(In229[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID230_INDEGREE3 n230 ( .InEdges(In230), .OutEdge(Out230),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID957 e957 ( .InEdge(Out134), .OutEdge(In230[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID958 e958 ( .InEdge(Out405), .OutEdge(In230[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID959 e959 ( .InEdge(Out387), .OutEdge(In230[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID231_INDEGREE3 n231 ( .InEdges(In231), .OutEdge(Out231),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID960 e960 ( .InEdge(Out278), .OutEdge(In231[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID961 e961 ( .InEdge(Out103), .OutEdge(In231[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID962 e962 ( .InEdge(Out379), .OutEdge(In231[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID232_INDEGREE1 n232 ( .InEdges(In232), .OutEdge(Out232),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID963 e963 ( .InEdge(Out311), .OutEdge(In232[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID233_INDEGREE6 n233 ( .InEdges(In233), .OutEdge(Out233),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID964 e964 ( .InEdge(Out314), .OutEdge(In233[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID965 e965 ( .InEdge(Out400), .OutEdge(In233[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID966 e966 ( .InEdge(Out161), .OutEdge(In233[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID967 e967 ( .InEdge(Out229), .OutEdge(In233[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID968 e968 ( .InEdge(Out406), .OutEdge(In233[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID969 e969 ( .InEdge(Out463), .OutEdge(In233[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID234_INDEGREE1 n234 ( .InEdges(In234), .OutEdge(Out234),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID970 e970 ( .InEdge(Out233), .OutEdge(In234[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID235_INDEGREE3 n235 ( .InEdges(In235), .OutEdge(Out235),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID971 e971 ( .InEdge(Out476), .OutEdge(In235[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID972 e972 ( .InEdge(Out218), .OutEdge(In235[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID973 e973 ( .InEdge(Out296), .OutEdge(In235[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID236_INDEGREE2 n236 ( .InEdges(In236), .OutEdge(Out236),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID974 e974 ( .InEdge(Out166), .OutEdge(In236[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID975 e975 ( .InEdge(Out380), .OutEdge(In236[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID237_INDEGREE4 n237 ( .InEdges(In237), .OutEdge(Out237),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID976 e976 ( .InEdge(Out26), .OutEdge(In237[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID977 e977 ( .InEdge(Out483), .OutEdge(In237[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID978 e978 ( .InEdge(Out101), .OutEdge(In237[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID979 e979 ( .InEdge(Out49), .OutEdge(In237[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID238_INDEGREE7 n238 ( .InEdges(In238), .OutEdge(Out238),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID980 e980 ( .InEdge(Out434), .OutEdge(In238[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID981 e981 ( .InEdge(Out436), .OutEdge(In238[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID982 e982 ( .InEdge(Out126), .OutEdge(In238[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID983 e983 ( .InEdge(Out237), .OutEdge(In238[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID984 e984 ( .InEdge(Out422), .OutEdge(In238[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID985 e985 ( .InEdge(Out210), .OutEdge(In238[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID986 e986 ( .InEdge(Out485), .OutEdge(In238[6:6]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID239_INDEGREE5 n239 ( .InEdges(In239), .OutEdge(Out239),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID987 e987 ( .InEdge(Out216), .OutEdge(In239[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID988 e988 ( .InEdge(Out420), .OutEdge(In239[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID989 e989 ( .InEdge(Out275), .OutEdge(In239[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID990 e990 ( .InEdge(Out212), .OutEdge(In239[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID991 e991 ( .InEdge(Out280), .OutEdge(In239[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID240_INDEGREE1 n240 ( .InEdges(In240), .OutEdge(Out240),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID992 e992 ( .InEdge(Out141), .OutEdge(In240[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID241_INDEGREE4 n241 ( .InEdges(In241), .OutEdge(Out241),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID993 e993 ( .InEdge(Out172), .OutEdge(In241[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID994 e994 ( .InEdge(Out168), .OutEdge(In241[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID995 e995 ( .InEdge(Out95), .OutEdge(In241[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID996 e996 ( .InEdge(Out509), .OutEdge(In241[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID242_INDEGREE4 n242 ( .InEdges(In242), .OutEdge(Out242),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID997 e997 ( .InEdge(Out389), .OutEdge(In242[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID998 e998 ( .InEdge(Out132), .OutEdge(In242[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID999 e999 ( .InEdge(Out158), .OutEdge(In242[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1000 e1000 ( .InEdge(Out137), .OutEdge(In242[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID243_INDEGREE3 n243 ( .InEdges(In243), .OutEdge(Out243),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1001 e1001 ( .InEdge(Out338), .OutEdge(In243[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1002 e1002 ( .InEdge(Out423), .OutEdge(In243[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1003 e1003 ( .InEdge(Out77), .OutEdge(In243[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID244_INDEGREE4 n244 ( .InEdges(In244), .OutEdge(Out244),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1004 e1004 ( .InEdge(Out407), .OutEdge(In244[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1005 e1005 ( .InEdge(Out253), .OutEdge(In244[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1006 e1006 ( .InEdge(Out156), .OutEdge(In244[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1007 e1007 ( .InEdge(Out452), .OutEdge(In244[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID245_INDEGREE3 n245 ( .InEdges(In245), .OutEdge(Out245),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1008 e1008 ( .InEdge(Out196), .OutEdge(In245[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1009 e1009 ( .InEdge(Out153), .OutEdge(In245[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1010 e1010 ( .InEdge(Out109), .OutEdge(In245[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID246_INDEGREE5 n246 ( .InEdges(In246), .OutEdge(Out246),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1011 e1011 ( .InEdge(Out158), .OutEdge(In246[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1012 e1012 ( .InEdge(Out181), .OutEdge(In246[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1013 e1013 ( .InEdge(Out353), .OutEdge(In246[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1014 e1014 ( .InEdge(Out446), .OutEdge(In246[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1015 e1015 ( .InEdge(Out178), .OutEdge(In246[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID247_INDEGREE5 n247 ( .InEdges(In247), .OutEdge(Out247),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1016 e1016 ( .InEdge(Out171), .OutEdge(In247[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1017 e1017 ( .InEdge(Out59), .OutEdge(In247[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1018 e1018 ( .InEdge(Out214), .OutEdge(In247[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1019 e1019 ( .InEdge(Out493), .OutEdge(In247[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1020 e1020 ( .InEdge(Out430), .OutEdge(In247[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID248_INDEGREE2 n248 ( .InEdges(In248), .OutEdge(Out248),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1021 e1021 ( .InEdge(Out410), .OutEdge(In248[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1022 e1022 ( .InEdge(Out77), .OutEdge(In248[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID249_INDEGREE7 n249 ( .InEdges(In249), .OutEdge(Out249),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1023 e1023 ( .InEdge(Out484), .OutEdge(In249[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1024 e1024 ( .InEdge(Out330), .OutEdge(In249[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1025 e1025 ( .InEdge(Out114), .OutEdge(In249[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1026 e1026 ( .InEdge(Out34), .OutEdge(In249[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1027 e1027 ( .InEdge(Out125), .OutEdge(In249[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1028 e1028 ( .InEdge(Out462), .OutEdge(In249[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1029 e1029 ( .InEdge(Out450), .OutEdge(In249[6:6]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID250_INDEGREE1 n250 ( .InEdges(In250), .OutEdge(Out250),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1030 e1030 ( .InEdge(Out140), .OutEdge(In250[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID251_INDEGREE5 n251 ( .InEdges(In251), .OutEdge(Out251),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1031 e1031 ( .InEdge(Out30), .OutEdge(In251[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1032 e1032 ( .InEdge(Out466), .OutEdge(In251[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1033 e1033 ( .InEdge(Out390), .OutEdge(In251[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1034 e1034 ( .InEdge(Out359), .OutEdge(In251[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1035 e1035 ( .InEdge(Out293), .OutEdge(In251[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID252_INDEGREE1 n252 ( .InEdges(In252), .OutEdge(Out252),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1036 e1036 ( .InEdge(Out454), .OutEdge(In252[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID253_INDEGREE2 n253 ( .InEdges(In253), .OutEdge(Out253),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1037 e1037 ( .InEdge(Out345), .OutEdge(In253[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1038 e1038 ( .InEdge(Out315), .OutEdge(In253[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID254_INDEGREE5 n254 ( .InEdges(In254), .OutEdge(Out254),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1039 e1039 ( .InEdge(Out491), .OutEdge(In254[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1040 e1040 ( .InEdge(Out379), .OutEdge(In254[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1041 e1041 ( .InEdge(Out351), .OutEdge(In254[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1042 e1042 ( .InEdge(Out54), .OutEdge(In254[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1043 e1043 ( .InEdge(Out431), .OutEdge(In254[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID255_INDEGREE1 n255 ( .InEdges(In255), .OutEdge(Out255),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1044 e1044 ( .InEdge(Out296), .OutEdge(In255[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID256_INDEGREE6 n256 ( .InEdges(In256), .OutEdge(Out256),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1045 e1045 ( .InEdge(Out65), .OutEdge(In256[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1046 e1046 ( .InEdge(Out66), .OutEdge(In256[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1047 e1047 ( .InEdge(Out477), .OutEdge(In256[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1048 e1048 ( .InEdge(Out496), .OutEdge(In256[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1049 e1049 ( .InEdge(Out313), .OutEdge(In256[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1050 e1050 ( .InEdge(Out271), .OutEdge(In256[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID257_INDEGREE3 n257 ( .InEdges(In257), .OutEdge(Out257),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1051 e1051 ( .InEdge(Out135), .OutEdge(In257[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1052 e1052 ( .InEdge(Out56), .OutEdge(In257[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1053 e1053 ( .InEdge(Out280), .OutEdge(In257[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID258_INDEGREE5 n258 ( .InEdges(In258), .OutEdge(Out258),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1054 e1054 ( .InEdge(Out403), .OutEdge(In258[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1055 e1055 ( .InEdge(Out143), .OutEdge(In258[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1056 e1056 ( .InEdge(Out310), .OutEdge(In258[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1057 e1057 ( .InEdge(Out396), .OutEdge(In258[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1058 e1058 ( .InEdge(Out364), .OutEdge(In258[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID259_INDEGREE4 n259 ( .InEdges(In259), .OutEdge(Out259),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1059 e1059 ( .InEdge(Out131), .OutEdge(In259[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1060 e1060 ( .InEdge(Out68), .OutEdge(In259[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1061 e1061 ( .InEdge(Out482), .OutEdge(In259[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1062 e1062 ( .InEdge(Out433), .OutEdge(In259[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID260_INDEGREE6 n260 ( .InEdges(In260), .OutEdge(Out260),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1063 e1063 ( .InEdge(Out352), .OutEdge(In260[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1064 e1064 ( .InEdge(Out402), .OutEdge(In260[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1065 e1065 ( .InEdge(Out284), .OutEdge(In260[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1066 e1066 ( .InEdge(Out280), .OutEdge(In260[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1067 e1067 ( .InEdge(Out187), .OutEdge(In260[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1068 e1068 ( .InEdge(Out105), .OutEdge(In260[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID261_INDEGREE3 n261 ( .InEdges(In261), .OutEdge(Out261),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1069 e1069 ( .InEdge(Out10), .OutEdge(In261[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1070 e1070 ( .InEdge(Out43), .OutEdge(In261[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1071 e1071 ( .InEdge(Out150), .OutEdge(In261[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID262_INDEGREE2 n262 ( .InEdges(In262), .OutEdge(Out262),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1072 e1072 ( .InEdge(Out209), .OutEdge(In262[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1073 e1073 ( .InEdge(Out79), .OutEdge(In262[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID263_INDEGREE3 n263 ( .InEdges(In263), .OutEdge(Out263),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1074 e1074 ( .InEdge(Out192), .OutEdge(In263[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1075 e1075 ( .InEdge(Out278), .OutEdge(In263[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1076 e1076 ( .InEdge(Out349), .OutEdge(In263[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID264_INDEGREE2 n264 ( .InEdges(In264), .OutEdge(Out264),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1077 e1077 ( .InEdge(Out128), .OutEdge(In264[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1078 e1078 ( .InEdge(Out74), .OutEdge(In264[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID265_INDEGREE1 n265 ( .InEdges(In265), .OutEdge(Out265),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1079 e1079 ( .InEdge(Out46), .OutEdge(In265[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID266_INDEGREE7 n266 ( .InEdges(In266), .OutEdge(Out266),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1080 e1080 ( .InEdge(Out189), .OutEdge(In266[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1081 e1081 ( .InEdge(Out123), .OutEdge(In266[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1082 e1082 ( .InEdge(Out312), .OutEdge(In266[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1083 e1083 ( .InEdge(Out218), .OutEdge(In266[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1084 e1084 ( .InEdge(Out37), .OutEdge(In266[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1085 e1085 ( .InEdge(Out8), .OutEdge(In266[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1086 e1086 ( .InEdge(Out416), .OutEdge(In266[6:6]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID267_INDEGREE5 n267 ( .InEdges(In267), .OutEdge(Out267),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1087 e1087 ( .InEdge(Out502), .OutEdge(In267[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1088 e1088 ( .InEdge(Out97), .OutEdge(In267[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1089 e1089 ( .InEdge(Out475), .OutEdge(In267[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1090 e1090 ( .InEdge(Out254), .OutEdge(In267[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1091 e1091 ( .InEdge(Out143), .OutEdge(In267[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID268_INDEGREE2 n268 ( .InEdges(In268), .OutEdge(Out268),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1092 e1092 ( .InEdge(Out301), .OutEdge(In268[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1093 e1093 ( .InEdge(Out401), .OutEdge(In268[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID269_INDEGREE1 n269 ( .InEdges(In269), .OutEdge(Out269),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1094 e1094 ( .InEdge(Out461), .OutEdge(In269[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID270_INDEGREE5 n270 ( .InEdges(In270), .OutEdge(Out270),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1095 e1095 ( .InEdge(Out402), .OutEdge(In270[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1096 e1096 ( .InEdge(Out174), .OutEdge(In270[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1097 e1097 ( .InEdge(Out186), .OutEdge(In270[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1098 e1098 ( .InEdge(Out114), .OutEdge(In270[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1099 e1099 ( .InEdge(Out92), .OutEdge(In270[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID271_INDEGREE5 n271 ( .InEdges(In271), .OutEdge(Out271),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1100 e1100 ( .InEdge(Out113), .OutEdge(In271[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1101 e1101 ( .InEdge(Out138), .OutEdge(In271[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1102 e1102 ( .InEdge(Out369), .OutEdge(In271[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1103 e1103 ( .InEdge(Out157), .OutEdge(In271[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1104 e1104 ( .InEdge(Out451), .OutEdge(In271[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID272_INDEGREE5 n272 ( .InEdges(In272), .OutEdge(Out272),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1105 e1105 ( .InEdge(Out369), .OutEdge(In272[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1106 e1106 ( .InEdge(Out497), .OutEdge(In272[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1107 e1107 ( .InEdge(Out261), .OutEdge(In272[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1108 e1108 ( .InEdge(Out273), .OutEdge(In272[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1109 e1109 ( .InEdge(Out306), .OutEdge(In272[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID273_INDEGREE7 n273 ( .InEdges(In273), .OutEdge(Out273),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1110 e1110 ( .InEdge(Out271), .OutEdge(In273[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1111 e1111 ( .InEdge(Out371), .OutEdge(In273[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1112 e1112 ( .InEdge(Out326), .OutEdge(In273[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1113 e1113 ( .InEdge(Out247), .OutEdge(In273[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1114 e1114 ( .InEdge(Out453), .OutEdge(In273[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1115 e1115 ( .InEdge(Out300), .OutEdge(In273[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1116 e1116 ( .InEdge(Out220), .OutEdge(In273[6:6]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID274_INDEGREE1 n274 ( .InEdges(In274), .OutEdge(Out274),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1117 e1117 ( .InEdge(Out451), .OutEdge(In274[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID275_INDEGREE1 n275 ( .InEdges(In275), .OutEdge(Out275),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1118 e1118 ( .InEdge(Out6), .OutEdge(In275[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID276_INDEGREE6 n276 ( .InEdges(In276), .OutEdge(Out276),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1119 e1119 ( .InEdge(Out511), .OutEdge(In276[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1120 e1120 ( .InEdge(Out368), .OutEdge(In276[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1121 e1121 ( .InEdge(Out403), .OutEdge(In276[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1122 e1122 ( .InEdge(Out391), .OutEdge(In276[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1123 e1123 ( .InEdge(Out72), .OutEdge(In276[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1124 e1124 ( .InEdge(Out396), .OutEdge(In276[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID277_INDEGREE1 n277 ( .InEdges(In277), .OutEdge(Out277),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1125 e1125 ( .InEdge(Out32), .OutEdge(In277[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID278_INDEGREE4 n278 ( .InEdges(In278), .OutEdge(Out278),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1126 e1126 ( .InEdge(Out193), .OutEdge(In278[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1127 e1127 ( .InEdge(Out186), .OutEdge(In278[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1128 e1128 ( .InEdge(Out367), .OutEdge(In278[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1129 e1129 ( .InEdge(Out314), .OutEdge(In278[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID279_INDEGREE1 n279 ( .InEdges(In279), .OutEdge(Out279),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1130 e1130 ( .InEdge(Out18), .OutEdge(In279[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID280_INDEGREE6 n280 ( .InEdges(In280), .OutEdge(Out280),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1131 e1131 ( .InEdge(Out66), .OutEdge(In280[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1132 e1132 ( .InEdge(Out179), .OutEdge(In280[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1133 e1133 ( .InEdge(Out362), .OutEdge(In280[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1134 e1134 ( .InEdge(Out506), .OutEdge(In280[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1135 e1135 ( .InEdge(Out208), .OutEdge(In280[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1136 e1136 ( .InEdge(Out339), .OutEdge(In280[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID281_INDEGREE3 n281 ( .InEdges(In281), .OutEdge(Out281),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1137 e1137 ( .InEdge(Out13), .OutEdge(In281[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1138 e1138 ( .InEdge(Out475), .OutEdge(In281[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1139 e1139 ( .InEdge(Out255), .OutEdge(In281[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID282_INDEGREE3 n282 ( .InEdges(In282), .OutEdge(Out282),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1140 e1140 ( .InEdge(Out394), .OutEdge(In282[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1141 e1141 ( .InEdge(Out355), .OutEdge(In282[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1142 e1142 ( .InEdge(Out431), .OutEdge(In282[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID283_INDEGREE7 n283 ( .InEdges(In283), .OutEdge(Out283),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1143 e1143 ( .InEdge(Out145), .OutEdge(In283[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1144 e1144 ( .InEdge(Out212), .OutEdge(In283[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1145 e1145 ( .InEdge(Out455), .OutEdge(In283[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1146 e1146 ( .InEdge(Out101), .OutEdge(In283[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1147 e1147 ( .InEdge(Out51), .OutEdge(In283[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1148 e1148 ( .InEdge(Out19), .OutEdge(In283[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1149 e1149 ( .InEdge(Out424), .OutEdge(In283[6:6]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID284_INDEGREE2 n284 ( .InEdges(In284), .OutEdge(Out284),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1150 e1150 ( .InEdge(Out281), .OutEdge(In284[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1151 e1151 ( .InEdge(Out408), .OutEdge(In284[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID285_INDEGREE2 n285 ( .InEdges(In285), .OutEdge(Out285),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1152 e1152 ( .InEdge(Out502), .OutEdge(In285[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1153 e1153 ( .InEdge(Out34), .OutEdge(In285[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID286_INDEGREE5 n286 ( .InEdges(In286), .OutEdge(Out286),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1154 e1154 ( .InEdge(Out14), .OutEdge(In286[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1155 e1155 ( .InEdge(Out143), .OutEdge(In286[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1156 e1156 ( .InEdge(Out182), .OutEdge(In286[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1157 e1157 ( .InEdge(Out277), .OutEdge(In286[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1158 e1158 ( .InEdge(Out407), .OutEdge(In286[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID287_INDEGREE1 n287 ( .InEdges(In287), .OutEdge(Out287),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1159 e1159 ( .InEdge(Out438), .OutEdge(In287[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID288_INDEGREE3 n288 ( .InEdges(In288), .OutEdge(Out288),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1160 e1160 ( .InEdge(Out398), .OutEdge(In288[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1161 e1161 ( .InEdge(Out480), .OutEdge(In288[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1162 e1162 ( .InEdge(Out488), .OutEdge(In288[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID289_INDEGREE2 n289 ( .InEdges(In289), .OutEdge(Out289),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1163 e1163 ( .InEdge(Out285), .OutEdge(In289[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1164 e1164 ( .InEdge(Out4), .OutEdge(In289[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID290_INDEGREE1 n290 ( .InEdges(In290), .OutEdge(Out290),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1165 e1165 ( .InEdge(Out336), .OutEdge(In290[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID291_INDEGREE3 n291 ( .InEdges(In291), .OutEdge(Out291),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1166 e1166 ( .InEdge(Out495), .OutEdge(In291[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1167 e1167 ( .InEdge(Out399), .OutEdge(In291[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1168 e1168 ( .InEdge(Out482), .OutEdge(In291[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID292_INDEGREE3 n292 ( .InEdges(In292), .OutEdge(Out292),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1169 e1169 ( .InEdge(Out500), .OutEdge(In292[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1170 e1170 ( .InEdge(Out138), .OutEdge(In292[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1171 e1171 ( .InEdge(Out195), .OutEdge(In292[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID293_INDEGREE1 n293 ( .InEdges(In293), .OutEdge(Out293),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1172 e1172 ( .InEdge(Out382), .OutEdge(In293[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID294_INDEGREE6 n294 ( .InEdges(In294), .OutEdge(Out294),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1173 e1173 ( .InEdge(Out216), .OutEdge(In294[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1174 e1174 ( .InEdge(Out398), .OutEdge(In294[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1175 e1175 ( .InEdge(Out481), .OutEdge(In294[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1176 e1176 ( .InEdge(Out417), .OutEdge(In294[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1177 e1177 ( .InEdge(Out151), .OutEdge(In294[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1178 e1178 ( .InEdge(Out466), .OutEdge(In294[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID295_INDEGREE5 n295 ( .InEdges(In295), .OutEdge(Out295),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1179 e1179 ( .InEdge(Out344), .OutEdge(In295[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1180 e1180 ( .InEdge(Out384), .OutEdge(In295[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1181 e1181 ( .InEdge(Out353), .OutEdge(In295[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1182 e1182 ( .InEdge(Out196), .OutEdge(In295[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1183 e1183 ( .InEdge(Out50), .OutEdge(In295[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID296_INDEGREE1 n296 ( .InEdges(In296), .OutEdge(Out296),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1184 e1184 ( .InEdge(Out68), .OutEdge(In296[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID297_INDEGREE5 n297 ( .InEdges(In297), .OutEdge(Out297),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1185 e1185 ( .InEdge(Out397), .OutEdge(In297[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1186 e1186 ( .InEdge(Out137), .OutEdge(In297[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1187 e1187 ( .InEdge(Out73), .OutEdge(In297[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1188 e1188 ( .InEdge(Out61), .OutEdge(In297[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1189 e1189 ( .InEdge(Out221), .OutEdge(In297[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID298_INDEGREE7 n298 ( .InEdges(In298), .OutEdge(Out298),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1190 e1190 ( .InEdge(Out102), .OutEdge(In298[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1191 e1191 ( .InEdge(Out301), .OutEdge(In298[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1192 e1192 ( .InEdge(Out203), .OutEdge(In298[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1193 e1193 ( .InEdge(Out464), .OutEdge(In298[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1194 e1194 ( .InEdge(Out384), .OutEdge(In298[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1195 e1195 ( .InEdge(Out483), .OutEdge(In298[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1196 e1196 ( .InEdge(Out34), .OutEdge(In298[6:6]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID299_INDEGREE7 n299 ( .InEdges(In299), .OutEdge(Out299),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1197 e1197 ( .InEdge(Out175), .OutEdge(In299[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1198 e1198 ( .InEdge(Out53), .OutEdge(In299[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1199 e1199 ( .InEdge(Out403), .OutEdge(In299[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1200 e1200 ( .InEdge(Out169), .OutEdge(In299[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1201 e1201 ( .InEdge(Out194), .OutEdge(In299[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1202 e1202 ( .InEdge(Out398), .OutEdge(In299[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1203 e1203 ( .InEdge(Out511), .OutEdge(In299[6:6]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID300_INDEGREE3 n300 ( .InEdges(In300), .OutEdge(Out300),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1204 e1204 ( .InEdge(Out273), .OutEdge(In300[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1205 e1205 ( .InEdge(Out283), .OutEdge(In300[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1206 e1206 ( .InEdge(Out271), .OutEdge(In300[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID301_INDEGREE2 n301 ( .InEdges(In301), .OutEdge(Out301),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1207 e1207 ( .InEdge(Out25), .OutEdge(In301[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1208 e1208 ( .InEdge(Out472), .OutEdge(In301[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID302_INDEGREE2 n302 ( .InEdges(In302), .OutEdge(Out302),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1209 e1209 ( .InEdge(Out364), .OutEdge(In302[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1210 e1210 ( .InEdge(Out142), .OutEdge(In302[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID303_INDEGREE7 n303 ( .InEdges(In303), .OutEdge(Out303),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1211 e1211 ( .InEdge(Out376), .OutEdge(In303[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1212 e1212 ( .InEdge(Out158), .OutEdge(In303[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1213 e1213 ( .InEdge(Out141), .OutEdge(In303[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1214 e1214 ( .InEdge(Out125), .OutEdge(In303[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1215 e1215 ( .InEdge(Out310), .OutEdge(In303[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1216 e1216 ( .InEdge(Out317), .OutEdge(In303[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1217 e1217 ( .InEdge(Out452), .OutEdge(In303[6:6]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID304_INDEGREE5 n304 ( .InEdges(In304), .OutEdge(Out304),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1218 e1218 ( .InEdge(Out410), .OutEdge(In304[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1219 e1219 ( .InEdge(Out361), .OutEdge(In304[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1220 e1220 ( .InEdge(Out367), .OutEdge(In304[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1221 e1221 ( .InEdge(Out13), .OutEdge(In304[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1222 e1222 ( .InEdge(Out510), .OutEdge(In304[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID305_INDEGREE3 n305 ( .InEdges(In305), .OutEdge(Out305),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1223 e1223 ( .InEdge(Out184), .OutEdge(In305[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1224 e1224 ( .InEdge(Out179), .OutEdge(In305[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1225 e1225 ( .InEdge(Out335), .OutEdge(In305[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID306_INDEGREE2 n306 ( .InEdges(In306), .OutEdge(Out306),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1226 e1226 ( .InEdge(Out327), .OutEdge(In306[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1227 e1227 ( .InEdge(Out97), .OutEdge(In306[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID307_INDEGREE2 n307 ( .InEdges(In307), .OutEdge(Out307),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1228 e1228 ( .InEdge(Out6), .OutEdge(In307[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1229 e1229 ( .InEdge(Out223), .OutEdge(In307[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID308_INDEGREE4 n308 ( .InEdges(In308), .OutEdge(Out308),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1230 e1230 ( .InEdge(Out443), .OutEdge(In308[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1231 e1231 ( .InEdge(Out141), .OutEdge(In308[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1232 e1232 ( .InEdge(Out109), .OutEdge(In308[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1233 e1233 ( .InEdge(Out377), .OutEdge(In308[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID309_INDEGREE5 n309 ( .InEdges(In309), .OutEdge(Out309),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1234 e1234 ( .InEdge(Out296), .OutEdge(In309[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1235 e1235 ( .InEdge(Out333), .OutEdge(In309[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1236 e1236 ( .InEdge(Out346), .OutEdge(In309[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1237 e1237 ( .InEdge(Out482), .OutEdge(In309[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1238 e1238 ( .InEdge(Out366), .OutEdge(In309[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID310_INDEGREE5 n310 ( .InEdges(In310), .OutEdge(Out310),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1239 e1239 ( .InEdge(Out113), .OutEdge(In310[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1240 e1240 ( .InEdge(Out353), .OutEdge(In310[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1241 e1241 ( .InEdge(Out10), .OutEdge(In310[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1242 e1242 ( .InEdge(Out222), .OutEdge(In310[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1243 e1243 ( .InEdge(Out308), .OutEdge(In310[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID311_INDEGREE4 n311 ( .InEdges(In311), .OutEdge(Out311),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1244 e1244 ( .InEdge(Out87), .OutEdge(In311[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1245 e1245 ( .InEdge(Out82), .OutEdge(In311[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1246 e1246 ( .InEdge(Out304), .OutEdge(In311[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1247 e1247 ( .InEdge(Out255), .OutEdge(In311[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID312_INDEGREE5 n312 ( .InEdges(In312), .OutEdge(Out312),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1248 e1248 ( .InEdge(Out351), .OutEdge(In312[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1249 e1249 ( .InEdge(Out253), .OutEdge(In312[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1250 e1250 ( .InEdge(Out6), .OutEdge(In312[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1251 e1251 ( .InEdge(Out493), .OutEdge(In312[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1252 e1252 ( .InEdge(Out15), .OutEdge(In312[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID313_INDEGREE2 n313 ( .InEdges(In313), .OutEdge(Out313),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1253 e1253 ( .InEdge(Out390), .OutEdge(In313[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1254 e1254 ( .InEdge(Out294), .OutEdge(In313[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID314_INDEGREE1 n314 ( .InEdges(In314), .OutEdge(Out314),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1255 e1255 ( .InEdge(Out289), .OutEdge(In314[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID315_INDEGREE6 n315 ( .InEdges(In315), .OutEdge(Out315),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1256 e1256 ( .InEdge(Out275), .OutEdge(In315[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1257 e1257 ( .InEdge(Out70), .OutEdge(In315[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1258 e1258 ( .InEdge(Out474), .OutEdge(In315[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1259 e1259 ( .InEdge(Out176), .OutEdge(In315[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1260 e1260 ( .InEdge(Out289), .OutEdge(In315[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1261 e1261 ( .InEdge(Out358), .OutEdge(In315[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID316_INDEGREE5 n316 ( .InEdges(In316), .OutEdge(Out316),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1262 e1262 ( .InEdge(Out80), .OutEdge(In316[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1263 e1263 ( .InEdge(Out392), .OutEdge(In316[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1264 e1264 ( .InEdge(Out439), .OutEdge(In316[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1265 e1265 ( .InEdge(Out238), .OutEdge(In316[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1266 e1266 ( .InEdge(Out6), .OutEdge(In316[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID317_INDEGREE4 n317 ( .InEdges(In317), .OutEdge(Out317),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1267 e1267 ( .InEdge(Out165), .OutEdge(In317[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1268 e1268 ( .InEdge(Out508), .OutEdge(In317[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1269 e1269 ( .InEdge(Out268), .OutEdge(In317[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1270 e1270 ( .InEdge(Out281), .OutEdge(In317[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID318_INDEGREE3 n318 ( .InEdges(In318), .OutEdge(Out318),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1271 e1271 ( .InEdge(Out493), .OutEdge(In318[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1272 e1272 ( .InEdge(Out76), .OutEdge(In318[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1273 e1273 ( .InEdge(Out144), .OutEdge(In318[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID319_INDEGREE1 n319 ( .InEdges(In319), .OutEdge(Out319),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1274 e1274 ( .InEdge(Out235), .OutEdge(In319[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID320_INDEGREE7 n320 ( .InEdges(In320), .OutEdge(Out320),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1275 e1275 ( .InEdge(Out507), .OutEdge(In320[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1276 e1276 ( .InEdge(Out440), .OutEdge(In320[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1277 e1277 ( .InEdge(Out421), .OutEdge(In320[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1278 e1278 ( .InEdge(Out315), .OutEdge(In320[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1279 e1279 ( .InEdge(Out112), .OutEdge(In320[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1280 e1280 ( .InEdge(Out16), .OutEdge(In320[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1281 e1281 ( .InEdge(Out230), .OutEdge(In320[6:6]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID321_INDEGREE1 n321 ( .InEdges(In321), .OutEdge(Out321),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1282 e1282 ( .InEdge(Out379), .OutEdge(In321[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID322_INDEGREE7 n322 ( .InEdges(In322), .OutEdge(Out322),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1283 e1283 ( .InEdge(Out52), .OutEdge(In322[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1284 e1284 ( .InEdge(Out366), .OutEdge(In322[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1285 e1285 ( .InEdge(Out472), .OutEdge(In322[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1286 e1286 ( .InEdge(Out167), .OutEdge(In322[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1287 e1287 ( .InEdge(Out362), .OutEdge(In322[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1288 e1288 ( .InEdge(Out356), .OutEdge(In322[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1289 e1289 ( .InEdge(Out41), .OutEdge(In322[6:6]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID323_INDEGREE3 n323 ( .InEdges(In323), .OutEdge(Out323),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1290 e1290 ( .InEdge(Out505), .OutEdge(In323[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1291 e1291 ( .InEdge(Out399), .OutEdge(In323[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1292 e1292 ( .InEdge(Out360), .OutEdge(In323[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID324_INDEGREE7 n324 ( .InEdges(In324), .OutEdge(Out324),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1293 e1293 ( .InEdge(Out474), .OutEdge(In324[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1294 e1294 ( .InEdge(Out138), .OutEdge(In324[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1295 e1295 ( .InEdge(Out145), .OutEdge(In324[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1296 e1296 ( .InEdge(Out285), .OutEdge(In324[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1297 e1297 ( .InEdge(Out238), .OutEdge(In324[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1298 e1298 ( .InEdge(Out290), .OutEdge(In324[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1299 e1299 ( .InEdge(Out209), .OutEdge(In324[6:6]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID325_INDEGREE2 n325 ( .InEdges(In325), .OutEdge(Out325),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1300 e1300 ( .InEdge(Out479), .OutEdge(In325[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1301 e1301 ( .InEdge(Out294), .OutEdge(In325[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID326_INDEGREE5 n326 ( .InEdges(In326), .OutEdge(Out326),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1302 e1302 ( .InEdge(Out342), .OutEdge(In326[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1303 e1303 ( .InEdge(Out202), .OutEdge(In326[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1304 e1304 ( .InEdge(Out314), .OutEdge(In326[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1305 e1305 ( .InEdge(Out79), .OutEdge(In326[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1306 e1306 ( .InEdge(Out222), .OutEdge(In326[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID327_INDEGREE3 n327 ( .InEdges(In327), .OutEdge(Out327),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1307 e1307 ( .InEdge(Out197), .OutEdge(In327[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1308 e1308 ( .InEdge(Out506), .OutEdge(In327[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1309 e1309 ( .InEdge(Out267), .OutEdge(In327[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID328_INDEGREE6 n328 ( .InEdges(In328), .OutEdge(Out328),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1310 e1310 ( .InEdge(Out45), .OutEdge(In328[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1311 e1311 ( .InEdge(Out110), .OutEdge(In328[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1312 e1312 ( .InEdge(Out293), .OutEdge(In328[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1313 e1313 ( .InEdge(Out359), .OutEdge(In328[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1314 e1314 ( .InEdge(Out415), .OutEdge(In328[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1315 e1315 ( .InEdge(Out62), .OutEdge(In328[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID329_INDEGREE7 n329 ( .InEdges(In329), .OutEdge(Out329),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1316 e1316 ( .InEdge(Out247), .OutEdge(In329[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1317 e1317 ( .InEdge(Out82), .OutEdge(In329[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1318 e1318 ( .InEdge(Out213), .OutEdge(In329[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1319 e1319 ( .InEdge(Out68), .OutEdge(In329[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1320 e1320 ( .InEdge(Out15), .OutEdge(In329[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1321 e1321 ( .InEdge(Out426), .OutEdge(In329[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1322 e1322 ( .InEdge(Out454), .OutEdge(In329[6:6]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID330_INDEGREE5 n330 ( .InEdges(In330), .OutEdge(Out330),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1323 e1323 ( .InEdge(Out38), .OutEdge(In330[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1324 e1324 ( .InEdge(Out101), .OutEdge(In330[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1325 e1325 ( .InEdge(Out277), .OutEdge(In330[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1326 e1326 ( .InEdge(Out336), .OutEdge(In330[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1327 e1327 ( .InEdge(Out359), .OutEdge(In330[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID331_INDEGREE6 n331 ( .InEdges(In331), .OutEdge(Out331),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1328 e1328 ( .InEdge(Out198), .OutEdge(In331[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1329 e1329 ( .InEdge(Out338), .OutEdge(In331[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1330 e1330 ( .InEdge(Out319), .OutEdge(In331[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1331 e1331 ( .InEdge(Out130), .OutEdge(In331[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1332 e1332 ( .InEdge(Out134), .OutEdge(In331[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1333 e1333 ( .InEdge(Out294), .OutEdge(In331[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID332_INDEGREE6 n332 ( .InEdges(In332), .OutEdge(Out332),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1334 e1334 ( .InEdge(Out301), .OutEdge(In332[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1335 e1335 ( .InEdge(Out504), .OutEdge(In332[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1336 e1336 ( .InEdge(Out135), .OutEdge(In332[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1337 e1337 ( .InEdge(Out57), .OutEdge(In332[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1338 e1338 ( .InEdge(Out65), .OutEdge(In332[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1339 e1339 ( .InEdge(Out495), .OutEdge(In332[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID333_INDEGREE4 n333 ( .InEdges(In333), .OutEdge(Out333),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1340 e1340 ( .InEdge(Out507), .OutEdge(In333[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1341 e1341 ( .InEdge(Out344), .OutEdge(In333[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1342 e1342 ( .InEdge(Out343), .OutEdge(In333[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1343 e1343 ( .InEdge(Out497), .OutEdge(In333[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID334_INDEGREE3 n334 ( .InEdges(In334), .OutEdge(Out334),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1344 e1344 ( .InEdge(Out300), .OutEdge(In334[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1345 e1345 ( .InEdge(Out371), .OutEdge(In334[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1346 e1346 ( .InEdge(Out356), .OutEdge(In334[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID335_INDEGREE5 n335 ( .InEdges(In335), .OutEdge(Out335),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1347 e1347 ( .InEdge(Out132), .OutEdge(In335[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1348 e1348 ( .InEdge(Out205), .OutEdge(In335[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1349 e1349 ( .InEdge(Out9), .OutEdge(In335[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1350 e1350 ( .InEdge(Out506), .OutEdge(In335[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1351 e1351 ( .InEdge(Out185), .OutEdge(In335[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID336_INDEGREE4 n336 ( .InEdges(In336), .OutEdge(Out336),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1352 e1352 ( .InEdge(Out289), .OutEdge(In336[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1353 e1353 ( .InEdge(Out324), .OutEdge(In336[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1354 e1354 ( .InEdge(Out426), .OutEdge(In336[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1355 e1355 ( .InEdge(Out123), .OutEdge(In336[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID337_INDEGREE3 n337 ( .InEdges(In337), .OutEdge(Out337),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1356 e1356 ( .InEdge(Out0), .OutEdge(In337[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1357 e1357 ( .InEdge(Out398), .OutEdge(In337[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1358 e1358 ( .InEdge(Out153), .OutEdge(In337[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID338_INDEGREE1 n338 ( .InEdges(In338), .OutEdge(Out338),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1359 e1359 ( .InEdge(Out466), .OutEdge(In338[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID339_INDEGREE3 n339 ( .InEdges(In339), .OutEdge(Out339),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1360 e1360 ( .InEdge(Out362), .OutEdge(In339[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1361 e1361 ( .InEdge(Out125), .OutEdge(In339[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1362 e1362 ( .InEdge(Out367), .OutEdge(In339[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID340_INDEGREE5 n340 ( .InEdges(In340), .OutEdge(Out340),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1363 e1363 ( .InEdge(Out491), .OutEdge(In340[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1364 e1364 ( .InEdge(Out374), .OutEdge(In340[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1365 e1365 ( .InEdge(Out472), .OutEdge(In340[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1366 e1366 ( .InEdge(Out209), .OutEdge(In340[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1367 e1367 ( .InEdge(Out107), .OutEdge(In340[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID341_INDEGREE6 n341 ( .InEdges(In341), .OutEdge(Out341),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1368 e1368 ( .InEdge(Out244), .OutEdge(In341[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1369 e1369 ( .InEdge(Out76), .OutEdge(In341[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1370 e1370 ( .InEdge(Out191), .OutEdge(In341[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1371 e1371 ( .InEdge(Out32), .OutEdge(In341[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1372 e1372 ( .InEdge(Out39), .OutEdge(In341[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1373 e1373 ( .InEdge(Out86), .OutEdge(In341[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID342_INDEGREE3 n342 ( .InEdges(In342), .OutEdge(Out342),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1374 e1374 ( .InEdge(Out387), .OutEdge(In342[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1375 e1375 ( .InEdge(Out402), .OutEdge(In342[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1376 e1376 ( .InEdge(Out18), .OutEdge(In342[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID343_INDEGREE1 n343 ( .InEdges(In343), .OutEdge(Out343),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1377 e1377 ( .InEdge(Out207), .OutEdge(In343[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID344_INDEGREE4 n344 ( .InEdges(In344), .OutEdge(Out344),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1378 e1378 ( .InEdge(Out429), .OutEdge(In344[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1379 e1379 ( .InEdge(Out306), .OutEdge(In344[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1380 e1380 ( .InEdge(Out40), .OutEdge(In344[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1381 e1381 ( .InEdge(Out451), .OutEdge(In344[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID345_INDEGREE5 n345 ( .InEdges(In345), .OutEdge(Out345),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1382 e1382 ( .InEdge(Out258), .OutEdge(In345[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1383 e1383 ( .InEdge(Out217), .OutEdge(In345[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1384 e1384 ( .InEdge(Out165), .OutEdge(In345[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1385 e1385 ( .InEdge(Out1), .OutEdge(In345[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1386 e1386 ( .InEdge(Out306), .OutEdge(In345[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID346_INDEGREE7 n346 ( .InEdges(In346), .OutEdge(Out346),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1387 e1387 ( .InEdge(Out94), .OutEdge(In346[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1388 e1388 ( .InEdge(Out244), .OutEdge(In346[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1389 e1389 ( .InEdge(Out261), .OutEdge(In346[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1390 e1390 ( .InEdge(Out131), .OutEdge(In346[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1391 e1391 ( .InEdge(Out66), .OutEdge(In346[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1392 e1392 ( .InEdge(Out9), .OutEdge(In346[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1393 e1393 ( .InEdge(Out103), .OutEdge(In346[6:6]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID347_INDEGREE3 n347 ( .InEdges(In347), .OutEdge(Out347),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1394 e1394 ( .InEdge(Out118), .OutEdge(In347[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1395 e1395 ( .InEdge(Out256), .OutEdge(In347[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1396 e1396 ( .InEdge(Out171), .OutEdge(In347[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID348_INDEGREE2 n348 ( .InEdges(In348), .OutEdge(Out348),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1397 e1397 ( .InEdge(Out173), .OutEdge(In348[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1398 e1398 ( .InEdge(Out457), .OutEdge(In348[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID349_INDEGREE2 n349 ( .InEdges(In349), .OutEdge(Out349),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1399 e1399 ( .InEdge(Out12), .OutEdge(In349[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1400 e1400 ( .InEdge(Out116), .OutEdge(In349[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID350_INDEGREE6 n350 ( .InEdges(In350), .OutEdge(Out350),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1401 e1401 ( .InEdge(Out17), .OutEdge(In350[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1402 e1402 ( .InEdge(Out48), .OutEdge(In350[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1403 e1403 ( .InEdge(Out437), .OutEdge(In350[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1404 e1404 ( .InEdge(Out418), .OutEdge(In350[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1405 e1405 ( .InEdge(Out454), .OutEdge(In350[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1406 e1406 ( .InEdge(Out478), .OutEdge(In350[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID351_INDEGREE2 n351 ( .InEdges(In351), .OutEdge(Out351),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1407 e1407 ( .InEdge(Out314), .OutEdge(In351[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1408 e1408 ( .InEdge(Out279), .OutEdge(In351[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID352_INDEGREE1 n352 ( .InEdges(In352), .OutEdge(Out352),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1409 e1409 ( .InEdge(Out401), .OutEdge(In352[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID353_INDEGREE4 n353 ( .InEdges(In353), .OutEdge(Out353),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1410 e1410 ( .InEdge(Out223), .OutEdge(In353[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1411 e1411 ( .InEdge(Out303), .OutEdge(In353[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1412 e1412 ( .InEdge(Out15), .OutEdge(In353[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1413 e1413 ( .InEdge(Out200), .OutEdge(In353[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID354_INDEGREE7 n354 ( .InEdges(In354), .OutEdge(Out354),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1414 e1414 ( .InEdge(Out311), .OutEdge(In354[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1415 e1415 ( .InEdge(Out3), .OutEdge(In354[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1416 e1416 ( .InEdge(Out352), .OutEdge(In354[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1417 e1417 ( .InEdge(Out406), .OutEdge(In354[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1418 e1418 ( .InEdge(Out380), .OutEdge(In354[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1419 e1419 ( .InEdge(Out501), .OutEdge(In354[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1420 e1420 ( .InEdge(Out254), .OutEdge(In354[6:6]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID355_INDEGREE4 n355 ( .InEdges(In355), .OutEdge(Out355),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1421 e1421 ( .InEdge(Out432), .OutEdge(In355[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1422 e1422 ( .InEdge(Out94), .OutEdge(In355[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1423 e1423 ( .InEdge(Out85), .OutEdge(In355[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1424 e1424 ( .InEdge(Out254), .OutEdge(In355[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID356_INDEGREE5 n356 ( .InEdges(In356), .OutEdge(Out356),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1425 e1425 ( .InEdge(Out23), .OutEdge(In356[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1426 e1426 ( .InEdge(Out259), .OutEdge(In356[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1427 e1427 ( .InEdge(Out442), .OutEdge(In356[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1428 e1428 ( .InEdge(Out458), .OutEdge(In356[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1429 e1429 ( .InEdge(Out257), .OutEdge(In356[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID357_INDEGREE1 n357 ( .InEdges(In357), .OutEdge(Out357),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1430 e1430 ( .InEdge(Out289), .OutEdge(In357[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID358_INDEGREE4 n358 ( .InEdges(In358), .OutEdge(Out358),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1431 e1431 ( .InEdge(Out51), .OutEdge(In358[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1432 e1432 ( .InEdge(Out230), .OutEdge(In358[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1433 e1433 ( .InEdge(Out164), .OutEdge(In358[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1434 e1434 ( .InEdge(Out356), .OutEdge(In358[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID359_INDEGREE6 n359 ( .InEdges(In359), .OutEdge(Out359),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1435 e1435 ( .InEdge(Out357), .OutEdge(In359[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1436 e1436 ( .InEdge(Out225), .OutEdge(In359[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1437 e1437 ( .InEdge(Out269), .OutEdge(In359[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1438 e1438 ( .InEdge(Out495), .OutEdge(In359[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1439 e1439 ( .InEdge(Out154), .OutEdge(In359[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1440 e1440 ( .InEdge(Out136), .OutEdge(In359[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID360_INDEGREE6 n360 ( .InEdges(In360), .OutEdge(Out360),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1441 e1441 ( .InEdge(Out215), .OutEdge(In360[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1442 e1442 ( .InEdge(Out90), .OutEdge(In360[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1443 e1443 ( .InEdge(Out153), .OutEdge(In360[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1444 e1444 ( .InEdge(Out274), .OutEdge(In360[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1445 e1445 ( .InEdge(Out5), .OutEdge(In360[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1446 e1446 ( .InEdge(Out365), .OutEdge(In360[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID361_INDEGREE5 n361 ( .InEdges(In361), .OutEdge(Out361),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1447 e1447 ( .InEdge(Out272), .OutEdge(In361[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1448 e1448 ( .InEdge(Out305), .OutEdge(In361[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1449 e1449 ( .InEdge(Out55), .OutEdge(In361[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1450 e1450 ( .InEdge(Out316), .OutEdge(In361[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1451 e1451 ( .InEdge(Out173), .OutEdge(In361[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID362_INDEGREE3 n362 ( .InEdges(In362), .OutEdge(Out362),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1452 e1452 ( .InEdge(Out232), .OutEdge(In362[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1453 e1453 ( .InEdge(Out340), .OutEdge(In362[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1454 e1454 ( .InEdge(Out282), .OutEdge(In362[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID363_INDEGREE3 n363 ( .InEdges(In363), .OutEdge(Out363),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1455 e1455 ( .InEdge(Out280), .OutEdge(In363[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1456 e1456 ( .InEdge(Out169), .OutEdge(In363[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1457 e1457 ( .InEdge(Out293), .OutEdge(In363[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID364_INDEGREE5 n364 ( .InEdges(In364), .OutEdge(Out364),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1458 e1458 ( .InEdge(Out160), .OutEdge(In364[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1459 e1459 ( .InEdge(Out452), .OutEdge(In364[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1460 e1460 ( .InEdge(Out196), .OutEdge(In364[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1461 e1461 ( .InEdge(Out314), .OutEdge(In364[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1462 e1462 ( .InEdge(Out13), .OutEdge(In364[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID365_INDEGREE3 n365 ( .InEdges(In365), .OutEdge(Out365),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1463 e1463 ( .InEdge(Out322), .OutEdge(In365[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1464 e1464 ( .InEdge(Out112), .OutEdge(In365[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1465 e1465 ( .InEdge(Out476), .OutEdge(In365[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID366_INDEGREE1 n366 ( .InEdges(In366), .OutEdge(Out366),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1466 e1466 ( .InEdge(Out216), .OutEdge(In366[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID367_INDEGREE6 n367 ( .InEdges(In367), .OutEdge(Out367),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1467 e1467 ( .InEdge(Out76), .OutEdge(In367[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1468 e1468 ( .InEdge(Out52), .OutEdge(In367[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1469 e1469 ( .InEdge(Out30), .OutEdge(In367[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1470 e1470 ( .InEdge(Out111), .OutEdge(In367[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1471 e1471 ( .InEdge(Out89), .OutEdge(In367[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1472 e1472 ( .InEdge(Out317), .OutEdge(In367[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID368_INDEGREE6 n368 ( .InEdges(In368), .OutEdge(Out368),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1473 e1473 ( .InEdge(Out132), .OutEdge(In368[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1474 e1474 ( .InEdge(Out399), .OutEdge(In368[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1475 e1475 ( .InEdge(Out225), .OutEdge(In368[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1476 e1476 ( .InEdge(Out115), .OutEdge(In368[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1477 e1477 ( .InEdge(Out141), .OutEdge(In368[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1478 e1478 ( .InEdge(Out164), .OutEdge(In368[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID369_INDEGREE5 n369 ( .InEdges(In369), .OutEdge(Out369),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1479 e1479 ( .InEdge(Out439), .OutEdge(In369[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1480 e1480 ( .InEdge(Out184), .OutEdge(In369[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1481 e1481 ( .InEdge(Out241), .OutEdge(In369[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1482 e1482 ( .InEdge(Out305), .OutEdge(In369[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1483 e1483 ( .InEdge(Out102), .OutEdge(In369[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID370_INDEGREE5 n370 ( .InEdges(In370), .OutEdge(Out370),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1484 e1484 ( .InEdge(Out479), .OutEdge(In370[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1485 e1485 ( .InEdge(Out292), .OutEdge(In370[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1486 e1486 ( .InEdge(Out146), .OutEdge(In370[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1487 e1487 ( .InEdge(Out53), .OutEdge(In370[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1488 e1488 ( .InEdge(Out15), .OutEdge(In370[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID371_INDEGREE7 n371 ( .InEdges(In371), .OutEdge(Out371),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1489 e1489 ( .InEdge(Out82), .OutEdge(In371[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1490 e1490 ( .InEdge(Out417), .OutEdge(In371[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1491 e1491 ( .InEdge(Out238), .OutEdge(In371[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1492 e1492 ( .InEdge(Out410), .OutEdge(In371[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1493 e1493 ( .InEdge(Out49), .OutEdge(In371[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1494 e1494 ( .InEdge(Out484), .OutEdge(In371[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1495 e1495 ( .InEdge(Out48), .OutEdge(In371[6:6]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID372_INDEGREE4 n372 ( .InEdges(In372), .OutEdge(Out372),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1496 e1496 ( .InEdge(Out467), .OutEdge(In372[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1497 e1497 ( .InEdge(Out280), .OutEdge(In372[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1498 e1498 ( .InEdge(Out140), .OutEdge(In372[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1499 e1499 ( .InEdge(Out479), .OutEdge(In372[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID373_INDEGREE2 n373 ( .InEdges(In373), .OutEdge(Out373),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1500 e1500 ( .InEdge(Out250), .OutEdge(In373[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1501 e1501 ( .InEdge(Out67), .OutEdge(In373[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID374_INDEGREE6 n374 ( .InEdges(In374), .OutEdge(Out374),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1502 e1502 ( .InEdge(Out413), .OutEdge(In374[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1503 e1503 ( .InEdge(Out52), .OutEdge(In374[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1504 e1504 ( .InEdge(Out109), .OutEdge(In374[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1505 e1505 ( .InEdge(Out329), .OutEdge(In374[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1506 e1506 ( .InEdge(Out225), .OutEdge(In374[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1507 e1507 ( .InEdge(Out389), .OutEdge(In374[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID375_INDEGREE2 n375 ( .InEdges(In375), .OutEdge(Out375),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1508 e1508 ( .InEdge(Out501), .OutEdge(In375[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1509 e1509 ( .InEdge(Out145), .OutEdge(In375[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID376_INDEGREE4 n376 ( .InEdges(In376), .OutEdge(Out376),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1510 e1510 ( .InEdge(Out285), .OutEdge(In376[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1511 e1511 ( .InEdge(Out370), .OutEdge(In376[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1512 e1512 ( .InEdge(Out23), .OutEdge(In376[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1513 e1513 ( .InEdge(Out310), .OutEdge(In376[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID377_INDEGREE4 n377 ( .InEdges(In377), .OutEdge(Out377),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1514 e1514 ( .InEdge(Out499), .OutEdge(In377[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1515 e1515 ( .InEdge(Out81), .OutEdge(In377[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1516 e1516 ( .InEdge(Out461), .OutEdge(In377[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1517 e1517 ( .InEdge(Out403), .OutEdge(In377[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID378_INDEGREE5 n378 ( .InEdges(In378), .OutEdge(Out378),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1518 e1518 ( .InEdge(Out119), .OutEdge(In378[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1519 e1519 ( .InEdge(Out309), .OutEdge(In378[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1520 e1520 ( .InEdge(Out45), .OutEdge(In378[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1521 e1521 ( .InEdge(Out25), .OutEdge(In378[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1522 e1522 ( .InEdge(Out465), .OutEdge(In378[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID379_INDEGREE4 n379 ( .InEdges(In379), .OutEdge(Out379),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1523 e1523 ( .InEdge(Out327), .OutEdge(In379[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1524 e1524 ( .InEdge(Out294), .OutEdge(In379[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1525 e1525 ( .InEdge(Out236), .OutEdge(In379[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1526 e1526 ( .InEdge(Out383), .OutEdge(In379[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID380_INDEGREE2 n380 ( .InEdges(In380), .OutEdge(Out380),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1527 e1527 ( .InEdge(Out205), .OutEdge(In380[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1528 e1528 ( .InEdge(Out208), .OutEdge(In380[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID381_INDEGREE5 n381 ( .InEdges(In381), .OutEdge(Out381),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1529 e1529 ( .InEdge(Out345), .OutEdge(In381[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1530 e1530 ( .InEdge(Out386), .OutEdge(In381[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1531 e1531 ( .InEdge(Out343), .OutEdge(In381[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1532 e1532 ( .InEdge(Out454), .OutEdge(In381[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1533 e1533 ( .InEdge(Out497), .OutEdge(In381[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID382_INDEGREE3 n382 ( .InEdges(In382), .OutEdge(Out382),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1534 e1534 ( .InEdge(Out453), .OutEdge(In382[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1535 e1535 ( .InEdge(Out182), .OutEdge(In382[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1536 e1536 ( .InEdge(Out243), .OutEdge(In382[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID383_INDEGREE3 n383 ( .InEdges(In383), .OutEdge(Out383),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1537 e1537 ( .InEdge(Out467), .OutEdge(In383[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1538 e1538 ( .InEdge(Out198), .OutEdge(In383[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1539 e1539 ( .InEdge(Out313), .OutEdge(In383[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID384_INDEGREE1 n384 ( .InEdges(In384), .OutEdge(Out384),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1540 e1540 ( .InEdge(Out410), .OutEdge(In384[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID385_INDEGREE3 n385 ( .InEdges(In385), .OutEdge(Out385),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1541 e1541 ( .InEdge(Out108), .OutEdge(In385[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1542 e1542 ( .InEdge(Out287), .OutEdge(In385[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1543 e1543 ( .InEdge(Out226), .OutEdge(In385[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID386_INDEGREE6 n386 ( .InEdges(In386), .OutEdge(Out386),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1544 e1544 ( .InEdge(Out68), .OutEdge(In386[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1545 e1545 ( .InEdge(Out355), .OutEdge(In386[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1546 e1546 ( .InEdge(Out434), .OutEdge(In386[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1547 e1547 ( .InEdge(Out128), .OutEdge(In386[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1548 e1548 ( .InEdge(Out232), .OutEdge(In386[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1549 e1549 ( .InEdge(Out17), .OutEdge(In386[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID387_INDEGREE7 n387 ( .InEdges(In387), .OutEdge(Out387),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1550 e1550 ( .InEdge(Out199), .OutEdge(In387[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1551 e1551 ( .InEdge(Out39), .OutEdge(In387[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1552 e1552 ( .InEdge(Out194), .OutEdge(In387[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1553 e1553 ( .InEdge(Out404), .OutEdge(In387[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1554 e1554 ( .InEdge(Out5), .OutEdge(In387[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1555 e1555 ( .InEdge(Out368), .OutEdge(In387[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1556 e1556 ( .InEdge(Out161), .OutEdge(In387[6:6]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID388_INDEGREE7 n388 ( .InEdges(In388), .OutEdge(Out388),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1557 e1557 ( .InEdge(Out122), .OutEdge(In388[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1558 e1558 ( .InEdge(Out155), .OutEdge(In388[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1559 e1559 ( .InEdge(Out164), .OutEdge(In388[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1560 e1560 ( .InEdge(Out57), .OutEdge(In388[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1561 e1561 ( .InEdge(Out127), .OutEdge(In388[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1562 e1562 ( .InEdge(Out470), .OutEdge(In388[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1563 e1563 ( .InEdge(Out431), .OutEdge(In388[6:6]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID389_INDEGREE4 n389 ( .InEdges(In389), .OutEdge(Out389),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1564 e1564 ( .InEdge(Out277), .OutEdge(In389[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1565 e1565 ( .InEdge(Out327), .OutEdge(In389[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1566 e1566 ( .InEdge(Out214), .OutEdge(In389[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1567 e1567 ( .InEdge(Out231), .OutEdge(In389[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID390_INDEGREE5 n390 ( .InEdges(In390), .OutEdge(Out390),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1568 e1568 ( .InEdge(Out482), .OutEdge(In390[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1569 e1569 ( .InEdge(Out194), .OutEdge(In390[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1570 e1570 ( .InEdge(Out38), .OutEdge(In390[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1571 e1571 ( .InEdge(Out438), .OutEdge(In390[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1572 e1572 ( .InEdge(Out195), .OutEdge(In390[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID391_INDEGREE6 n391 ( .InEdges(In391), .OutEdge(Out391),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1573 e1573 ( .InEdge(Out34), .OutEdge(In391[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1574 e1574 ( .InEdge(Out322), .OutEdge(In391[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1575 e1575 ( .InEdge(Out453), .OutEdge(In391[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1576 e1576 ( .InEdge(Out408), .OutEdge(In391[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1577 e1577 ( .InEdge(Out175), .OutEdge(In391[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1578 e1578 ( .InEdge(Out247), .OutEdge(In391[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID392_INDEGREE5 n392 ( .InEdges(In392), .OutEdge(Out392),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1579 e1579 ( .InEdge(Out342), .OutEdge(In392[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1580 e1580 ( .InEdge(Out149), .OutEdge(In392[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1581 e1581 ( .InEdge(Out462), .OutEdge(In392[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1582 e1582 ( .InEdge(Out331), .OutEdge(In392[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1583 e1583 ( .InEdge(Out485), .OutEdge(In392[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID393_INDEGREE6 n393 ( .InEdges(In393), .OutEdge(Out393),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1584 e1584 ( .InEdge(Out80), .OutEdge(In393[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1585 e1585 ( .InEdge(Out198), .OutEdge(In393[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1586 e1586 ( .InEdge(Out42), .OutEdge(In393[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1587 e1587 ( .InEdge(Out483), .OutEdge(In393[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1588 e1588 ( .InEdge(Out72), .OutEdge(In393[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1589 e1589 ( .InEdge(Out352), .OutEdge(In393[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID394_INDEGREE1 n394 ( .InEdges(In394), .OutEdge(Out394),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1590 e1590 ( .InEdge(Out476), .OutEdge(In394[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID395_INDEGREE1 n395 ( .InEdges(In395), .OutEdge(Out395),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1591 e1591 ( .InEdge(Out62), .OutEdge(In395[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID396_INDEGREE7 n396 ( .InEdges(In396), .OutEdge(Out396),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1592 e1592 ( .InEdge(Out480), .OutEdge(In396[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1593 e1593 ( .InEdge(Out122), .OutEdge(In396[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1594 e1594 ( .InEdge(Out121), .OutEdge(In396[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1595 e1595 ( .InEdge(Out510), .OutEdge(In396[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1596 e1596 ( .InEdge(Out415), .OutEdge(In396[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1597 e1597 ( .InEdge(Out11), .OutEdge(In396[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1598 e1598 ( .InEdge(Out412), .OutEdge(In396[6:6]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID397_INDEGREE6 n397 ( .InEdges(In397), .OutEdge(Out397),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1599 e1599 ( .InEdge(Out0), .OutEdge(In397[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1600 e1600 ( .InEdge(Out464), .OutEdge(In397[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1601 e1601 ( .InEdge(Out367), .OutEdge(In397[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1602 e1602 ( .InEdge(Out219), .OutEdge(In397[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1603 e1603 ( .InEdge(Out109), .OutEdge(In397[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1604 e1604 ( .InEdge(Out320), .OutEdge(In397[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID398_INDEGREE4 n398 ( .InEdges(In398), .OutEdge(Out398),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1605 e1605 ( .InEdge(Out383), .OutEdge(In398[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1606 e1606 ( .InEdge(Out438), .OutEdge(In398[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1607 e1607 ( .InEdge(Out347), .OutEdge(In398[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1608 e1608 ( .InEdge(Out337), .OutEdge(In398[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID399_INDEGREE5 n399 ( .InEdges(In399), .OutEdge(Out399),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1609 e1609 ( .InEdge(Out225), .OutEdge(In399[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1610 e1610 ( .InEdge(Out295), .OutEdge(In399[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1611 e1611 ( .InEdge(Out329), .OutEdge(In399[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1612 e1612 ( .InEdge(Out298), .OutEdge(In399[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1613 e1613 ( .InEdge(Out147), .OutEdge(In399[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID400_INDEGREE7 n400 ( .InEdges(In400), .OutEdge(Out400),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1614 e1614 ( .InEdge(Out107), .OutEdge(In400[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1615 e1615 ( .InEdge(Out385), .OutEdge(In400[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1616 e1616 ( .InEdge(Out77), .OutEdge(In400[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1617 e1617 ( .InEdge(Out8), .OutEdge(In400[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1618 e1618 ( .InEdge(Out451), .OutEdge(In400[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1619 e1619 ( .InEdge(Out484), .OutEdge(In400[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1620 e1620 ( .InEdge(Out392), .OutEdge(In400[6:6]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID401_INDEGREE7 n401 ( .InEdges(In401), .OutEdge(Out401),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1621 e1621 ( .InEdge(Out240), .OutEdge(In401[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1622 e1622 ( .InEdge(Out452), .OutEdge(In401[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1623 e1623 ( .InEdge(Out355), .OutEdge(In401[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1624 e1624 ( .InEdge(Out41), .OutEdge(In401[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1625 e1625 ( .InEdge(Out183), .OutEdge(In401[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1626 e1626 ( .InEdge(Out184), .OutEdge(In401[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1627 e1627 ( .InEdge(Out51), .OutEdge(In401[6:6]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID402_INDEGREE7 n402 ( .InEdges(In402), .OutEdge(Out402),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1628 e1628 ( .InEdge(Out496), .OutEdge(In402[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1629 e1629 ( .InEdge(Out327), .OutEdge(In402[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1630 e1630 ( .InEdge(Out108), .OutEdge(In402[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1631 e1631 ( .InEdge(Out481), .OutEdge(In402[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1632 e1632 ( .InEdge(Out410), .OutEdge(In402[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1633 e1633 ( .InEdge(Out210), .OutEdge(In402[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1634 e1634 ( .InEdge(Out3), .OutEdge(In402[6:6]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID403_INDEGREE7 n403 ( .InEdges(In403), .OutEdge(Out403),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1635 e1635 ( .InEdge(Out400), .OutEdge(In403[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1636 e1636 ( .InEdge(Out459), .OutEdge(In403[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1637 e1637 ( .InEdge(Out455), .OutEdge(In403[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1638 e1638 ( .InEdge(Out398), .OutEdge(In403[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1639 e1639 ( .InEdge(Out303), .OutEdge(In403[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1640 e1640 ( .InEdge(Out503), .OutEdge(In403[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1641 e1641 ( .InEdge(Out115), .OutEdge(In403[6:6]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID404_INDEGREE2 n404 ( .InEdges(In404), .OutEdge(Out404),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1642 e1642 ( .InEdge(Out408), .OutEdge(In404[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1643 e1643 ( .InEdge(Out88), .OutEdge(In404[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID405_INDEGREE6 n405 ( .InEdges(In405), .OutEdge(Out405),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1644 e1644 ( .InEdge(Out77), .OutEdge(In405[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1645 e1645 ( .InEdge(Out452), .OutEdge(In405[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1646 e1646 ( .InEdge(Out340), .OutEdge(In405[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1647 e1647 ( .InEdge(Out42), .OutEdge(In405[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1648 e1648 ( .InEdge(Out173), .OutEdge(In405[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1649 e1649 ( .InEdge(Out150), .OutEdge(In405[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID406_INDEGREE1 n406 ( .InEdges(In406), .OutEdge(Out406),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1650 e1650 ( .InEdge(Out47), .OutEdge(In406[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID407_INDEGREE2 n407 ( .InEdges(In407), .OutEdge(Out407),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1651 e1651 ( .InEdge(Out130), .OutEdge(In407[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1652 e1652 ( .InEdge(Out468), .OutEdge(In407[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID408_INDEGREE6 n408 ( .InEdges(In408), .OutEdge(Out408),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1653 e1653 ( .InEdge(Out221), .OutEdge(In408[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1654 e1654 ( .InEdge(Out328), .OutEdge(In408[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1655 e1655 ( .InEdge(Out13), .OutEdge(In408[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1656 e1656 ( .InEdge(Out220), .OutEdge(In408[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1657 e1657 ( .InEdge(Out49), .OutEdge(In408[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1658 e1658 ( .InEdge(Out381), .OutEdge(In408[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID409_INDEGREE4 n409 ( .InEdges(In409), .OutEdge(Out409),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1659 e1659 ( .InEdge(Out241), .OutEdge(In409[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1660 e1660 ( .InEdge(Out242), .OutEdge(In409[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1661 e1661 ( .InEdge(Out428), .OutEdge(In409[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1662 e1662 ( .InEdge(Out133), .OutEdge(In409[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID410_INDEGREE2 n410 ( .InEdges(In410), .OutEdge(Out410),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1663 e1663 ( .InEdge(Out496), .OutEdge(In410[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1664 e1664 ( .InEdge(Out316), .OutEdge(In410[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID411_INDEGREE1 n411 ( .InEdges(In411), .OutEdge(Out411),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1665 e1665 ( .InEdge(Out335), .OutEdge(In411[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID412_INDEGREE4 n412 ( .InEdges(In412), .OutEdge(Out412),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1666 e1666 ( .InEdge(Out401), .OutEdge(In412[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1667 e1667 ( .InEdge(Out42), .OutEdge(In412[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1668 e1668 ( .InEdge(Out491), .OutEdge(In412[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1669 e1669 ( .InEdge(Out107), .OutEdge(In412[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID413_INDEGREE4 n413 ( .InEdges(In413), .OutEdge(Out413),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1670 e1670 ( .InEdge(Out61), .OutEdge(In413[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1671 e1671 ( .InEdge(Out434), .OutEdge(In413[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1672 e1672 ( .InEdge(Out94), .OutEdge(In413[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1673 e1673 ( .InEdge(Out219), .OutEdge(In413[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID414_INDEGREE7 n414 ( .InEdges(In414), .OutEdge(Out414),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1674 e1674 ( .InEdge(Out324), .OutEdge(In414[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1675 e1675 ( .InEdge(Out43), .OutEdge(In414[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1676 e1676 ( .InEdge(Out63), .OutEdge(In414[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1677 e1677 ( .InEdge(Out510), .OutEdge(In414[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1678 e1678 ( .InEdge(Out34), .OutEdge(In414[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1679 e1679 ( .InEdge(Out360), .OutEdge(In414[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1680 e1680 ( .InEdge(Out480), .OutEdge(In414[6:6]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID415_INDEGREE4 n415 ( .InEdges(In415), .OutEdge(Out415),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1681 e1681 ( .InEdge(Out156), .OutEdge(In415[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1682 e1682 ( .InEdge(Out367), .OutEdge(In415[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1683 e1683 ( .InEdge(Out467), .OutEdge(In415[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1684 e1684 ( .InEdge(Out280), .OutEdge(In415[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID416_INDEGREE5 n416 ( .InEdges(In416), .OutEdge(Out416),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1685 e1685 ( .InEdge(Out486), .OutEdge(In416[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1686 e1686 ( .InEdge(Out255), .OutEdge(In416[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1687 e1687 ( .InEdge(Out163), .OutEdge(In416[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1688 e1688 ( .InEdge(Out348), .OutEdge(In416[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1689 e1689 ( .InEdge(Out466), .OutEdge(In416[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID417_INDEGREE3 n417 ( .InEdges(In417), .OutEdge(Out417),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1690 e1690 ( .InEdge(Out428), .OutEdge(In417[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1691 e1691 ( .InEdge(Out227), .OutEdge(In417[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1692 e1692 ( .InEdge(Out2), .OutEdge(In417[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID418_INDEGREE3 n418 ( .InEdges(In418), .OutEdge(Out418),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1693 e1693 ( .InEdge(Out473), .OutEdge(In418[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1694 e1694 ( .InEdge(Out137), .OutEdge(In418[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1695 e1695 ( .InEdge(Out290), .OutEdge(In418[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID419_INDEGREE6 n419 ( .InEdges(In419), .OutEdge(Out419),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1696 e1696 ( .InEdge(Out208), .OutEdge(In419[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1697 e1697 ( .InEdge(Out184), .OutEdge(In419[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1698 e1698 ( .InEdge(Out356), .OutEdge(In419[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1699 e1699 ( .InEdge(Out325), .OutEdge(In419[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1700 e1700 ( .InEdge(Out221), .OutEdge(In419[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1701 e1701 ( .InEdge(Out10), .OutEdge(In419[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID420_INDEGREE2 n420 ( .InEdges(In420), .OutEdge(Out420),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1702 e1702 ( .InEdge(Out190), .OutEdge(In420[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1703 e1703 ( .InEdge(Out150), .OutEdge(In420[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID421_INDEGREE6 n421 ( .InEdges(In421), .OutEdge(Out421),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1704 e1704 ( .InEdge(Out370), .OutEdge(In421[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1705 e1705 ( .InEdge(Out411), .OutEdge(In421[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1706 e1706 ( .InEdge(Out27), .OutEdge(In421[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1707 e1707 ( .InEdge(Out53), .OutEdge(In421[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1708 e1708 ( .InEdge(Out307), .OutEdge(In421[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1709 e1709 ( .InEdge(Out337), .OutEdge(In421[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID422_INDEGREE3 n422 ( .InEdges(In422), .OutEdge(Out422),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1710 e1710 ( .InEdge(Out483), .OutEdge(In422[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1711 e1711 ( .InEdge(Out317), .OutEdge(In422[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1712 e1712 ( .InEdge(Out157), .OutEdge(In422[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID423_INDEGREE1 n423 ( .InEdges(In423), .OutEdge(Out423),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1713 e1713 ( .InEdge(Out103), .OutEdge(In423[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID424_INDEGREE6 n424 ( .InEdges(In424), .OutEdge(Out424),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1714 e1714 ( .InEdge(Out410), .OutEdge(In424[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1715 e1715 ( .InEdge(Out248), .OutEdge(In424[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1716 e1716 ( .InEdge(Out147), .OutEdge(In424[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1717 e1717 ( .InEdge(Out278), .OutEdge(In424[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1718 e1718 ( .InEdge(Out405), .OutEdge(In424[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1719 e1719 ( .InEdge(Out374), .OutEdge(In424[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID425_INDEGREE2 n425 ( .InEdges(In425), .OutEdge(Out425),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1720 e1720 ( .InEdge(Out8), .OutEdge(In425[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1721 e1721 ( .InEdge(Out64), .OutEdge(In425[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID426_INDEGREE7 n426 ( .InEdges(In426), .OutEdge(Out426),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1722 e1722 ( .InEdge(Out102), .OutEdge(In426[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1723 e1723 ( .InEdge(Out393), .OutEdge(In426[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1724 e1724 ( .InEdge(Out361), .OutEdge(In426[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1725 e1725 ( .InEdge(Out157), .OutEdge(In426[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1726 e1726 ( .InEdge(Out278), .OutEdge(In426[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1727 e1727 ( .InEdge(Out248), .OutEdge(In426[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1728 e1728 ( .InEdge(Out178), .OutEdge(In426[6:6]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID427_INDEGREE1 n427 ( .InEdges(In427), .OutEdge(Out427),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1729 e1729 ( .InEdge(Out436), .OutEdge(In427[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID428_INDEGREE2 n428 ( .InEdges(In428), .OutEdge(Out428),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1730 e1730 ( .InEdge(Out416), .OutEdge(In428[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1731 e1731 ( .InEdge(Out457), .OutEdge(In428[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID429_INDEGREE1 n429 ( .InEdges(In429), .OutEdge(Out429),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1732 e1732 ( .InEdge(Out180), .OutEdge(In429[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID430_INDEGREE1 n430 ( .InEdges(In430), .OutEdge(Out430),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1733 e1733 ( .InEdge(Out110), .OutEdge(In430[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID431_INDEGREE1 n431 ( .InEdges(In431), .OutEdge(Out431),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1734 e1734 ( .InEdge(Out51), .OutEdge(In431[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID432_INDEGREE3 n432 ( .InEdges(In432), .OutEdge(Out432),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1735 e1735 ( .InEdge(Out380), .OutEdge(In432[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1736 e1736 ( .InEdge(Out30), .OutEdge(In432[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1737 e1737 ( .InEdge(Out331), .OutEdge(In432[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID433_INDEGREE7 n433 ( .InEdges(In433), .OutEdge(Out433),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1738 e1738 ( .InEdge(Out509), .OutEdge(In433[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1739 e1739 ( .InEdge(Out374), .OutEdge(In433[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1740 e1740 ( .InEdge(Out383), .OutEdge(In433[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1741 e1741 ( .InEdge(Out191), .OutEdge(In433[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1742 e1742 ( .InEdge(Out391), .OutEdge(In433[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1743 e1743 ( .InEdge(Out475), .OutEdge(In433[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1744 e1744 ( .InEdge(Out149), .OutEdge(In433[6:6]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID434_INDEGREE6 n434 ( .InEdges(In434), .OutEdge(Out434),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1745 e1745 ( .InEdge(Out43), .OutEdge(In434[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1746 e1746 ( .InEdge(Out143), .OutEdge(In434[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1747 e1747 ( .InEdge(Out203), .OutEdge(In434[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1748 e1748 ( .InEdge(Out354), .OutEdge(In434[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1749 e1749 ( .InEdge(Out209), .OutEdge(In434[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1750 e1750 ( .InEdge(Out80), .OutEdge(In434[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID435_INDEGREE2 n435 ( .InEdges(In435), .OutEdge(Out435),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1751 e1751 ( .InEdge(Out166), .OutEdge(In435[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1752 e1752 ( .InEdge(Out228), .OutEdge(In435[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID436_INDEGREE7 n436 ( .InEdges(In436), .OutEdge(Out436),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1753 e1753 ( .InEdge(Out457), .OutEdge(In436[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1754 e1754 ( .InEdge(Out217), .OutEdge(In436[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1755 e1755 ( .InEdge(Out388), .OutEdge(In436[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1756 e1756 ( .InEdge(Out151), .OutEdge(In436[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1757 e1757 ( .InEdge(Out280), .OutEdge(In436[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1758 e1758 ( .InEdge(Out264), .OutEdge(In436[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1759 e1759 ( .InEdge(Out362), .OutEdge(In436[6:6]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID437_INDEGREE4 n437 ( .InEdges(In437), .OutEdge(Out437),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1760 e1760 ( .InEdge(Out289), .OutEdge(In437[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1761 e1761 ( .InEdge(Out307), .OutEdge(In437[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1762 e1762 ( .InEdge(Out74), .OutEdge(In437[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1763 e1763 ( .InEdge(Out96), .OutEdge(In437[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID438_INDEGREE3 n438 ( .InEdges(In438), .OutEdge(Out438),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1764 e1764 ( .InEdge(Out117), .OutEdge(In438[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1765 e1765 ( .InEdge(Out122), .OutEdge(In438[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1766 e1766 ( .InEdge(Out368), .OutEdge(In438[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID439_INDEGREE1 n439 ( .InEdges(In439), .OutEdge(Out439),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1767 e1767 ( .InEdge(Out135), .OutEdge(In439[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID440_INDEGREE7 n440 ( .InEdges(In440), .OutEdge(Out440),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1768 e1768 ( .InEdge(Out288), .OutEdge(In440[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1769 e1769 ( .InEdge(Out125), .OutEdge(In440[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1770 e1770 ( .InEdge(Out0), .OutEdge(In440[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1771 e1771 ( .InEdge(Out484), .OutEdge(In440[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1772 e1772 ( .InEdge(Out403), .OutEdge(In440[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1773 e1773 ( .InEdge(Out309), .OutEdge(In440[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1774 e1774 ( .InEdge(Out425), .OutEdge(In440[6:6]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID441_INDEGREE3 n441 ( .InEdges(In441), .OutEdge(Out441),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1775 e1775 ( .InEdge(Out320), .OutEdge(In441[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1776 e1776 ( .InEdge(Out336), .OutEdge(In441[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1777 e1777 ( .InEdge(Out500), .OutEdge(In441[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID442_INDEGREE2 n442 ( .InEdges(In442), .OutEdge(Out442),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1778 e1778 ( .InEdge(Out0), .OutEdge(In442[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1779 e1779 ( .InEdge(Out430), .OutEdge(In442[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID443_INDEGREE6 n443 ( .InEdges(In443), .OutEdge(Out443),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1780 e1780 ( .InEdge(Out173), .OutEdge(In443[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1781 e1781 ( .InEdge(Out482), .OutEdge(In443[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1782 e1782 ( .InEdge(Out270), .OutEdge(In443[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1783 e1783 ( .InEdge(Out334), .OutEdge(In443[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1784 e1784 ( .InEdge(Out502), .OutEdge(In443[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1785 e1785 ( .InEdge(Out392), .OutEdge(In443[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID444_INDEGREE2 n444 ( .InEdges(In444), .OutEdge(Out444),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1786 e1786 ( .InEdge(Out344), .OutEdge(In444[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1787 e1787 ( .InEdge(Out207), .OutEdge(In444[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID445_INDEGREE3 n445 ( .InEdges(In445), .OutEdge(Out445),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1788 e1788 ( .InEdge(Out109), .OutEdge(In445[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1789 e1789 ( .InEdge(Out500), .OutEdge(In445[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1790 e1790 ( .InEdge(Out354), .OutEdge(In445[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID446_INDEGREE4 n446 ( .InEdges(In446), .OutEdge(Out446),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1791 e1791 ( .InEdge(Out183), .OutEdge(In446[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1792 e1792 ( .InEdge(Out198), .OutEdge(In446[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1793 e1793 ( .InEdge(Out160), .OutEdge(In446[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1794 e1794 ( .InEdge(Out346), .OutEdge(In446[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID447_INDEGREE1 n447 ( .InEdges(In447), .OutEdge(Out447),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1795 e1795 ( .InEdge(Out385), .OutEdge(In447[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID448_INDEGREE3 n448 ( .InEdges(In448), .OutEdge(Out448),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1796 e1796 ( .InEdge(Out79), .OutEdge(In448[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1797 e1797 ( .InEdge(Out193), .OutEdge(In448[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1798 e1798 ( .InEdge(Out107), .OutEdge(In448[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID449_INDEGREE7 n449 ( .InEdges(In449), .OutEdge(Out449),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1799 e1799 ( .InEdge(Out452), .OutEdge(In449[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1800 e1800 ( .InEdge(Out32), .OutEdge(In449[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1801 e1801 ( .InEdge(Out232), .OutEdge(In449[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1802 e1802 ( .InEdge(Out354), .OutEdge(In449[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1803 e1803 ( .InEdge(Out338), .OutEdge(In449[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1804 e1804 ( .InEdge(Out504), .OutEdge(In449[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1805 e1805 ( .InEdge(Out195), .OutEdge(In449[6:6]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID450_INDEGREE4 n450 ( .InEdges(In450), .OutEdge(Out450),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1806 e1806 ( .InEdge(Out353), .OutEdge(In450[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1807 e1807 ( .InEdge(Out497), .OutEdge(In450[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1808 e1808 ( .InEdge(Out148), .OutEdge(In450[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1809 e1809 ( .InEdge(Out278), .OutEdge(In450[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID451_INDEGREE1 n451 ( .InEdges(In451), .OutEdge(Out451),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1810 e1810 ( .InEdge(Out143), .OutEdge(In451[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID452_INDEGREE2 n452 ( .InEdges(In452), .OutEdge(Out452),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1811 e1811 ( .InEdge(Out251), .OutEdge(In452[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1812 e1812 ( .InEdge(Out78), .OutEdge(In452[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID453_INDEGREE5 n453 ( .InEdges(In453), .OutEdge(Out453),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1813 e1813 ( .InEdge(Out368), .OutEdge(In453[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1814 e1814 ( .InEdge(Out31), .OutEdge(In453[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1815 e1815 ( .InEdge(Out394), .OutEdge(In453[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1816 e1816 ( .InEdge(Out118), .OutEdge(In453[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1817 e1817 ( .InEdge(Out295), .OutEdge(In453[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID454_INDEGREE5 n454 ( .InEdges(In454), .OutEdge(Out454),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1818 e1818 ( .InEdge(Out314), .OutEdge(In454[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1819 e1819 ( .InEdge(Out86), .OutEdge(In454[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1820 e1820 ( .InEdge(Out279), .OutEdge(In454[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1821 e1821 ( .InEdge(Out362), .OutEdge(In454[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1822 e1822 ( .InEdge(Out125), .OutEdge(In454[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID455_INDEGREE7 n455 ( .InEdges(In455), .OutEdge(Out455),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1823 e1823 ( .InEdge(Out39), .OutEdge(In455[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1824 e1824 ( .InEdge(Out191), .OutEdge(In455[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1825 e1825 ( .InEdge(Out30), .OutEdge(In455[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1826 e1826 ( .InEdge(Out62), .OutEdge(In455[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1827 e1827 ( .InEdge(Out422), .OutEdge(In455[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1828 e1828 ( .InEdge(Out167), .OutEdge(In455[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1829 e1829 ( .InEdge(Out306), .OutEdge(In455[6:6]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID456_INDEGREE2 n456 ( .InEdges(In456), .OutEdge(Out456),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1830 e1830 ( .InEdge(Out56), .OutEdge(In456[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1831 e1831 ( .InEdge(Out278), .OutEdge(In456[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID457_INDEGREE6 n457 ( .InEdges(In457), .OutEdge(Out457),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1832 e1832 ( .InEdge(Out23), .OutEdge(In457[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1833 e1833 ( .InEdge(Out312), .OutEdge(In457[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1834 e1834 ( .InEdge(Out161), .OutEdge(In457[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1835 e1835 ( .InEdge(Out57), .OutEdge(In457[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1836 e1836 ( .InEdge(Out110), .OutEdge(In457[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1837 e1837 ( .InEdge(Out355), .OutEdge(In457[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID458_INDEGREE7 n458 ( .InEdges(In458), .OutEdge(Out458),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1838 e1838 ( .InEdge(Out135), .OutEdge(In458[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1839 e1839 ( .InEdge(Out252), .OutEdge(In458[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1840 e1840 ( .InEdge(Out171), .OutEdge(In458[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1841 e1841 ( .InEdge(Out130), .OutEdge(In458[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1842 e1842 ( .InEdge(Out459), .OutEdge(In458[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1843 e1843 ( .InEdge(Out165), .OutEdge(In458[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1844 e1844 ( .InEdge(Out413), .OutEdge(In458[6:6]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID459_INDEGREE5 n459 ( .InEdges(In459), .OutEdge(Out459),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1845 e1845 ( .InEdge(Out380), .OutEdge(In459[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1846 e1846 ( .InEdge(Out375), .OutEdge(In459[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1847 e1847 ( .InEdge(Out184), .OutEdge(In459[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1848 e1848 ( .InEdge(Out150), .OutEdge(In459[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1849 e1849 ( .InEdge(Out170), .OutEdge(In459[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID460_INDEGREE7 n460 ( .InEdges(In460), .OutEdge(Out460),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1850 e1850 ( .InEdge(Out73), .OutEdge(In460[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1851 e1851 ( .InEdge(Out347), .OutEdge(In460[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1852 e1852 ( .InEdge(Out190), .OutEdge(In460[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1853 e1853 ( .InEdge(Out258), .OutEdge(In460[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1854 e1854 ( .InEdge(Out69), .OutEdge(In460[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1855 e1855 ( .InEdge(Out404), .OutEdge(In460[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1856 e1856 ( .InEdge(Out303), .OutEdge(In460[6:6]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID461_INDEGREE1 n461 ( .InEdges(In461), .OutEdge(Out461),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1857 e1857 ( .InEdge(Out355), .OutEdge(In461[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID462_INDEGREE6 n462 ( .InEdges(In462), .OutEdge(Out462),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1858 e1858 ( .InEdge(Out99), .OutEdge(In462[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1859 e1859 ( .InEdge(Out257), .OutEdge(In462[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1860 e1860 ( .InEdge(Out301), .OutEdge(In462[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1861 e1861 ( .InEdge(Out215), .OutEdge(In462[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1862 e1862 ( .InEdge(Out134), .OutEdge(In462[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1863 e1863 ( .InEdge(Out401), .OutEdge(In462[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID463_INDEGREE1 n463 ( .InEdges(In463), .OutEdge(Out463),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1864 e1864 ( .InEdge(Out271), .OutEdge(In463[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID464_INDEGREE4 n464 ( .InEdges(In464), .OutEdge(Out464),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1865 e1865 ( .InEdge(Out461), .OutEdge(In464[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1866 e1866 ( .InEdge(Out169), .OutEdge(In464[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1867 e1867 ( .InEdge(Out336), .OutEdge(In464[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1868 e1868 ( .InEdge(Out130), .OutEdge(In464[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID465_INDEGREE7 n465 ( .InEdges(In465), .OutEdge(Out465),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1869 e1869 ( .InEdge(Out240), .OutEdge(In465[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1870 e1870 ( .InEdge(Out277), .OutEdge(In465[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1871 e1871 ( .InEdge(Out116), .OutEdge(In465[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1872 e1872 ( .InEdge(Out12), .OutEdge(In465[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1873 e1873 ( .InEdge(Out392), .OutEdge(In465[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1874 e1874 ( .InEdge(Out86), .OutEdge(In465[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1875 e1875 ( .InEdge(Out345), .OutEdge(In465[6:6]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID466_INDEGREE4 n466 ( .InEdges(In466), .OutEdge(Out466),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1876 e1876 ( .InEdge(Out193), .OutEdge(In466[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1877 e1877 ( .InEdge(Out443), .OutEdge(In466[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1878 e1878 ( .InEdge(Out135), .OutEdge(In466[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1879 e1879 ( .InEdge(Out298), .OutEdge(In466[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID467_INDEGREE5 n467 ( .InEdges(In467), .OutEdge(Out467),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1880 e1880 ( .InEdge(Out204), .OutEdge(In467[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1881 e1881 ( .InEdge(Out101), .OutEdge(In467[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1882 e1882 ( .InEdge(Out452), .OutEdge(In467[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1883 e1883 ( .InEdge(Out432), .OutEdge(In467[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1884 e1884 ( .InEdge(Out234), .OutEdge(In467[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID468_INDEGREE1 n468 ( .InEdges(In468), .OutEdge(Out468),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1885 e1885 ( .InEdge(Out289), .OutEdge(In468[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID469_INDEGREE4 n469 ( .InEdges(In469), .OutEdge(Out469),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1886 e1886 ( .InEdge(Out6), .OutEdge(In469[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1887 e1887 ( .InEdge(Out430), .OutEdge(In469[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1888 e1888 ( .InEdge(Out414), .OutEdge(In469[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1889 e1889 ( .InEdge(Out242), .OutEdge(In469[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID470_INDEGREE2 n470 ( .InEdges(In470), .OutEdge(Out470),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1890 e1890 ( .InEdge(Out430), .OutEdge(In470[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1891 e1891 ( .InEdge(Out216), .OutEdge(In470[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID471_INDEGREE4 n471 ( .InEdges(In471), .OutEdge(Out471),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1892 e1892 ( .InEdge(Out508), .OutEdge(In471[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1893 e1893 ( .InEdge(Out160), .OutEdge(In471[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1894 e1894 ( .InEdge(Out11), .OutEdge(In471[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1895 e1895 ( .InEdge(Out414), .OutEdge(In471[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID472_INDEGREE6 n472 ( .InEdges(In472), .OutEdge(Out472),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1896 e1896 ( .InEdge(Out508), .OutEdge(In472[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1897 e1897 ( .InEdge(Out279), .OutEdge(In472[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1898 e1898 ( .InEdge(Out345), .OutEdge(In472[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1899 e1899 ( .InEdge(Out299), .OutEdge(In472[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1900 e1900 ( .InEdge(Out316), .OutEdge(In472[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1901 e1901 ( .InEdge(Out6), .OutEdge(In472[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID473_INDEGREE2 n473 ( .InEdges(In473), .OutEdge(Out473),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1902 e1902 ( .InEdge(Out175), .OutEdge(In473[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1903 e1903 ( .InEdge(Out287), .OutEdge(In473[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID474_INDEGREE2 n474 ( .InEdges(In474), .OutEdge(Out474),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1904 e1904 ( .InEdge(Out328), .OutEdge(In474[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1905 e1905 ( .InEdge(Out163), .OutEdge(In474[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID475_INDEGREE7 n475 ( .InEdges(In475), .OutEdge(Out475),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1906 e1906 ( .InEdge(Out266), .OutEdge(In475[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1907 e1907 ( .InEdge(Out325), .OutEdge(In475[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1908 e1908 ( .InEdge(Out105), .OutEdge(In475[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1909 e1909 ( .InEdge(Out409), .OutEdge(In475[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1910 e1910 ( .InEdge(Out51), .OutEdge(In475[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1911 e1911 ( .InEdge(Out214), .OutEdge(In475[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1912 e1912 ( .InEdge(Out164), .OutEdge(In475[6:6]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID476_INDEGREE5 n476 ( .InEdges(In476), .OutEdge(Out476),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1913 e1913 ( .InEdge(Out129), .OutEdge(In476[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1914 e1914 ( .InEdge(Out333), .OutEdge(In476[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1915 e1915 ( .InEdge(Out334), .OutEdge(In476[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1916 e1916 ( .InEdge(Out331), .OutEdge(In476[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1917 e1917 ( .InEdge(Out398), .OutEdge(In476[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID477_INDEGREE1 n477 ( .InEdges(In477), .OutEdge(Out477),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1918 e1918 ( .InEdge(Out106), .OutEdge(In477[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID478_INDEGREE7 n478 ( .InEdges(In478), .OutEdge(Out478),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1919 e1919 ( .InEdge(Out258), .OutEdge(In478[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1920 e1920 ( .InEdge(Out341), .OutEdge(In478[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1921 e1921 ( .InEdge(Out157), .OutEdge(In478[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1922 e1922 ( .InEdge(Out75), .OutEdge(In478[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1923 e1923 ( .InEdge(Out172), .OutEdge(In478[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1924 e1924 ( .InEdge(Out316), .OutEdge(In478[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1925 e1925 ( .InEdge(Out363), .OutEdge(In478[6:6]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID479_INDEGREE4 n479 ( .InEdges(In479), .OutEdge(Out479),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1926 e1926 ( .InEdge(Out502), .OutEdge(In479[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1927 e1927 ( .InEdge(Out266), .OutEdge(In479[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1928 e1928 ( .InEdge(Out103), .OutEdge(In479[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1929 e1929 ( .InEdge(Out390), .OutEdge(In479[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID480_INDEGREE5 n480 ( .InEdges(In480), .OutEdge(Out480),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1930 e1930 ( .InEdge(Out10), .OutEdge(In480[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1931 e1931 ( .InEdge(Out268), .OutEdge(In480[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1932 e1932 ( .InEdge(Out19), .OutEdge(In480[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1933 e1933 ( .InEdge(Out328), .OutEdge(In480[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1934 e1934 ( .InEdge(Out291), .OutEdge(In480[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID481_INDEGREE2 n481 ( .InEdges(In481), .OutEdge(Out481),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1935 e1935 ( .InEdge(Out201), .OutEdge(In481[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1936 e1936 ( .InEdge(Out372), .OutEdge(In481[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID482_INDEGREE3 n482 ( .InEdges(In482), .OutEdge(Out482),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1937 e1937 ( .InEdge(Out510), .OutEdge(In482[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1938 e1938 ( .InEdge(Out475), .OutEdge(In482[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1939 e1939 ( .InEdge(Out502), .OutEdge(In482[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID483_INDEGREE3 n483 ( .InEdges(In483), .OutEdge(Out483),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1940 e1940 ( .InEdge(Out379), .OutEdge(In483[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1941 e1941 ( .InEdge(Out343), .OutEdge(In483[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1942 e1942 ( .InEdge(Out106), .OutEdge(In483[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID484_INDEGREE2 n484 ( .InEdges(In484), .OutEdge(Out484),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1943 e1943 ( .InEdge(Out325), .OutEdge(In484[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1944 e1944 ( .InEdge(Out409), .OutEdge(In484[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID485_INDEGREE1 n485 ( .InEdges(In485), .OutEdge(Out485),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1945 e1945 ( .InEdge(Out319), .OutEdge(In485[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID486_INDEGREE1 n486 ( .InEdges(In486), .OutEdge(Out486),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1946 e1946 ( .InEdge(Out482), .OutEdge(In486[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID487_INDEGREE1 n487 ( .InEdges(In487), .OutEdge(Out487),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1947 e1947 ( .InEdge(Out274), .OutEdge(In487[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID488_INDEGREE7 n488 ( .InEdges(In488), .OutEdge(Out488),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1948 e1948 ( .InEdge(Out353), .OutEdge(In488[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1949 e1949 ( .InEdge(Out210), .OutEdge(In488[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1950 e1950 ( .InEdge(Out24), .OutEdge(In488[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1951 e1951 ( .InEdge(Out276), .OutEdge(In488[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1952 e1952 ( .InEdge(Out362), .OutEdge(In488[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1953 e1953 ( .InEdge(Out510), .OutEdge(In488[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1954 e1954 ( .InEdge(Out260), .OutEdge(In488[6:6]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID489_INDEGREE2 n489 ( .InEdges(In489), .OutEdge(Out489),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1955 e1955 ( .InEdge(Out111), .OutEdge(In489[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1956 e1956 ( .InEdge(Out28), .OutEdge(In489[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID490_INDEGREE4 n490 ( .InEdges(In490), .OutEdge(Out490),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1957 e1957 ( .InEdge(Out365), .OutEdge(In490[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1958 e1958 ( .InEdge(Out320), .OutEdge(In490[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1959 e1959 ( .InEdge(Out265), .OutEdge(In490[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1960 e1960 ( .InEdge(Out379), .OutEdge(In490[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID491_INDEGREE3 n491 ( .InEdges(In491), .OutEdge(Out491),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1961 e1961 ( .InEdge(Out318), .OutEdge(In491[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1962 e1962 ( .InEdge(Out89), .OutEdge(In491[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1963 e1963 ( .InEdge(Out74), .OutEdge(In491[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID492_INDEGREE5 n492 ( .InEdges(In492), .OutEdge(Out492),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1964 e1964 ( .InEdge(Out256), .OutEdge(In492[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1965 e1965 ( .InEdge(Out337), .OutEdge(In492[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1966 e1966 ( .InEdge(Out341), .OutEdge(In492[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1967 e1967 ( .InEdge(Out280), .OutEdge(In492[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1968 e1968 ( .InEdge(Out191), .OutEdge(In492[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID493_INDEGREE7 n493 ( .InEdges(In493), .OutEdge(Out493),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1969 e1969 ( .InEdge(Out32), .OutEdge(In493[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1970 e1970 ( .InEdge(Out356), .OutEdge(In493[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1971 e1971 ( .InEdge(Out390), .OutEdge(In493[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1972 e1972 ( .InEdge(Out258), .OutEdge(In493[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1973 e1973 ( .InEdge(Out238), .OutEdge(In493[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1974 e1974 ( .InEdge(Out257), .OutEdge(In493[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1975 e1975 ( .InEdge(Out108), .OutEdge(In493[6:6]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID494_INDEGREE3 n494 ( .InEdges(In494), .OutEdge(Out494),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1976 e1976 ( .InEdge(Out132), .OutEdge(In494[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1977 e1977 ( .InEdge(Out29), .OutEdge(In494[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1978 e1978 ( .InEdge(Out421), .OutEdge(In494[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID495_INDEGREE3 n495 ( .InEdges(In495), .OutEdge(Out495),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1979 e1979 ( .InEdge(Out81), .OutEdge(In495[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1980 e1980 ( .InEdge(Out274), .OutEdge(In495[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1981 e1981 ( .InEdge(Out332), .OutEdge(In495[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID496_INDEGREE4 n496 ( .InEdges(In496), .OutEdge(Out496),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1982 e1982 ( .InEdge(Out402), .OutEdge(In496[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1983 e1983 ( .InEdge(Out129), .OutEdge(In496[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1984 e1984 ( .InEdge(Out31), .OutEdge(In496[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1985 e1985 ( .InEdge(Out273), .OutEdge(In496[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID497_INDEGREE6 n497 ( .InEdges(In497), .OutEdge(Out497),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1986 e1986 ( .InEdge(Out16), .OutEdge(In497[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1987 e1987 ( .InEdge(Out463), .OutEdge(In497[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1988 e1988 ( .InEdge(Out400), .OutEdge(In497[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1989 e1989 ( .InEdge(Out386), .OutEdge(In497[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1990 e1990 ( .InEdge(Out250), .OutEdge(In497[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1991 e1991 ( .InEdge(Out410), .OutEdge(In497[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID498_INDEGREE5 n498 ( .InEdges(In498), .OutEdge(Out498),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1992 e1992 ( .InEdge(Out174), .OutEdge(In498[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1993 e1993 ( .InEdge(Out467), .OutEdge(In498[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1994 e1994 ( .InEdge(Out462), .OutEdge(In498[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1995 e1995 ( .InEdge(Out420), .OutEdge(In498[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1996 e1996 ( .InEdge(Out71), .OutEdge(In498[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID499_INDEGREE4 n499 ( .InEdges(In499), .OutEdge(Out499),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID1997 e1997 ( .InEdge(Out385), .OutEdge(In499[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1998 e1998 ( .InEdge(Out207), .OutEdge(In499[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID1999 e1999 ( .InEdge(Out81), .OutEdge(In499[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID2000 e2000 ( .InEdge(Out333), .OutEdge(In499[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID500_INDEGREE1 n500 ( .InEdges(In500), .OutEdge(Out500),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID2001 e2001 ( .InEdge(Out245), .OutEdge(In500[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID501_INDEGREE4 n501 ( .InEdges(In501), .OutEdge(Out501),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID2002 e2002 ( .InEdge(Out470), .OutEdge(In501[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID2003 e2003 ( .InEdge(Out255), .OutEdge(In501[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID2004 e2004 ( .InEdge(Out370), .OutEdge(In501[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID2005 e2005 ( .InEdge(Out216), .OutEdge(In501[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID502_INDEGREE6 n502 ( .InEdges(In502), .OutEdge(Out502),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID2006 e2006 ( .InEdge(Out108), .OutEdge(In502[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID2007 e2007 ( .InEdge(Out347), .OutEdge(In502[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID2008 e2008 ( .InEdge(Out134), .OutEdge(In502[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID2009 e2009 ( .InEdge(Out358), .OutEdge(In502[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID2010 e2010 ( .InEdge(Out118), .OutEdge(In502[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID2011 e2011 ( .InEdge(Out310), .OutEdge(In502[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID503_INDEGREE7 n503 ( .InEdges(In503), .OutEdge(Out503),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID2012 e2012 ( .InEdge(Out463), .OutEdge(In503[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID2013 e2013 ( .InEdge(Out63), .OutEdge(In503[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID2014 e2014 ( .InEdge(Out134), .OutEdge(In503[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID2015 e2015 ( .InEdge(Out61), .OutEdge(In503[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID2016 e2016 ( .InEdge(Out446), .OutEdge(In503[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID2017 e2017 ( .InEdge(Out57), .OutEdge(In503[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID2018 e2018 ( .InEdge(Out158), .OutEdge(In503[6:6]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID504_INDEGREE1 n504 ( .InEdges(In504), .OutEdge(Out504),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID2019 e2019 ( .InEdge(Out46), .OutEdge(In504[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID505_INDEGREE7 n505 ( .InEdges(In505), .OutEdge(Out505),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID2020 e2020 ( .InEdge(Out72), .OutEdge(In505[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID2021 e2021 ( .InEdge(Out417), .OutEdge(In505[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID2022 e2022 ( .InEdge(Out180), .OutEdge(In505[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID2023 e2023 ( .InEdge(Out273), .OutEdge(In505[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID2024 e2024 ( .InEdge(Out82), .OutEdge(In505[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID2025 e2025 ( .InEdge(Out492), .OutEdge(In505[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID2026 e2026 ( .InEdge(Out449), .OutEdge(In505[6:6]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID506_INDEGREE6 n506 ( .InEdges(In506), .OutEdge(Out506),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID2027 e2027 ( .InEdge(Out94), .OutEdge(In506[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID2028 e2028 ( .InEdge(Out78), .OutEdge(In506[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID2029 e2029 ( .InEdge(Out421), .OutEdge(In506[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID2030 e2030 ( .InEdge(Out361), .OutEdge(In506[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID2031 e2031 ( .InEdge(Out389), .OutEdge(In506[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID2032 e2032 ( .InEdge(Out68), .OutEdge(In506[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID507_INDEGREE5 n507 ( .InEdges(In507), .OutEdge(Out507),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID2033 e2033 ( .InEdge(Out90), .OutEdge(In507[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID2034 e2034 ( .InEdge(Out32), .OutEdge(In507[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID2035 e2035 ( .InEdge(Out130), .OutEdge(In507[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID2036 e2036 ( .InEdge(Out466), .OutEdge(In507[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID2037 e2037 ( .InEdge(Out456), .OutEdge(In507[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID508_INDEGREE7 n508 ( .InEdges(In508), .OutEdge(Out508),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID2038 e2038 ( .InEdge(Out17), .OutEdge(In508[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID2039 e2039 ( .InEdge(Out343), .OutEdge(In508[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID2040 e2040 ( .InEdge(Out270), .OutEdge(In508[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID2041 e2041 ( .InEdge(Out436), .OutEdge(In508[3:3]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID2042 e2042 ( .InEdge(Out305), .OutEdge(In508[4:4]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID2043 e2043 ( .InEdge(Out494), .OutEdge(In508[5:5]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID2044 e2044 ( .InEdge(Out287), .OutEdge(In508[6:6]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID509_INDEGREE1 n509 ( .InEdges(In509), .OutEdge(Out509),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID2045 e2045 ( .InEdge(Out237), .OutEdge(In509[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID510_INDEGREE3 n510 ( .InEdges(In510), .OutEdge(Out510),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID2046 e2046 ( .InEdge(Out443), .OutEdge(In510[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID2047 e2047 ( .InEdge(Out429), .OutEdge(In510[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID2048 e2048 ( .InEdge(Out480), .OutEdge(In510[2:2]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );

    Node_NID511_INDEGREE2 n511 ( .InEdges(In511), .OutEdge(Out511),
        .PathAddr(PathAddr), .PathData(PathData),
        .Start(Start), .Clk(Clk) );
    Edge_EID2049 e2049 ( .InEdge(Out2), .OutEdge(In511[0:0]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
    Edge_EID2050 e2050 ( .InEdge(Out502), .OutEdge(In511[1:1]),
        .WeightAddr(WeightAddr), .WeightData(WeightData),
        .Clk(Clk) );
endmodule
